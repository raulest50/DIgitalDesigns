-- megafunction wizard: %ALTFP_SINCOS%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altfp_sincos 

-- ============================================================
-- File Name: mysincos.vhd
-- Megafunction Name(s):
-- 			altfp_sincos
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altfp_sincos CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" OPERATION="SIN" PIPELINE=36 ROUNDING="TO_NEAREST" WIDTH_EXP=8 WIDTH_MAN=23 clock data result
--VERSION_BEGIN 13.0 cbx_altfp_sincos 2013:06:12:18:03:43:SJ cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_clshift 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END


--altfp_sincos_cordic_m CBX_AUTO_BLACKBOX="ALL" DEPTH=18 DEVICE_FAMILY="Cyclone II" INDEXPOINT=2 WIDTH=34 aclr clken clock indexbit radians sincos sincosbit
--VERSION_BEGIN 13.0 cbx_altfp_sincos 2013:06:12:18:03:43:SJ cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_clshift 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" indexpoint=2 START=0 WIDTH=34 arctan indexbit
--VERSION_BEGIN 13.0 cbx_altfp_sincos 2013:06:12:18:03:43:SJ cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_clshift 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altfp_sincos_cordic_atan_08b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END mysincos_altfp_sincos_cordic_atan_08b;

 ARCHITECTURE RTL OF mysincos_altfp_sincos_cordic_atan_08b IS

	 SIGNAL  wire_cata_0_cordic_atan_w_lg_w_lg_indexbit10924w10925w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_0_cordic_atan_w_lg_indexbit10922w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_0_cordic_atan_w_lg_indexbit10924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_0_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_2_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_0_cordic_atan_w_valuenode_0_w_range10923w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_0_cordic_atan_w_valuenode_2_w_range10921w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop0 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_0_cordic_atan_w_lg_w_lg_indexbit10924w10925w(i) <= wire_cata_0_cordic_atan_w_lg_indexbit10924w(0) AND wire_cata_0_cordic_atan_w_valuenode_0_w_range10923w(i);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_0_cordic_atan_w_lg_indexbit10922w(i) <= indexbit AND wire_cata_0_cordic_atan_w_valuenode_2_w_range10921w(i);
	END GENERATE loop1;
	wire_cata_0_cordic_atan_w_lg_indexbit10924w(0) <= NOT indexbit;
	arctan <= (wire_cata_0_cordic_atan_w_lg_w_lg_indexbit10924w10925w OR wire_cata_0_cordic_atan_w_lg_indexbit10922w);
	valuenode_0_w <= "001100100100001111110110101010001000100001011010";
	valuenode_2_w <= "000011111010110110111010111111001001011001000000";
	wire_cata_0_cordic_atan_w_valuenode_0_w_range10923w <= valuenode_0_w(47 DOWNTO 14);
	wire_cata_0_cordic_atan_w_valuenode_2_w_range10921w <= valuenode_2_w(45 DOWNTO 12);

 END RTL; --mysincos_altfp_sincos_cordic_atan_08b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" indexpoint=2 START=10 WIDTH=34 arctan indexbit
--VERSION_BEGIN 13.0 cbx_altfp_sincos 2013:06:12:18:03:43:SJ cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_clshift 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altfp_sincos_cordic_atan_h9b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END mysincos_altfp_sincos_cordic_atan_h9b;

 ARCHITECTURE RTL OF mysincos_altfp_sincos_cordic_atan_h9b IS

	 SIGNAL  wire_cata_10_cordic_atan_w_lg_w_lg_indexbit10930w10931w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_10_cordic_atan_w_lg_indexbit10928w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_10_cordic_atan_w_lg_indexbit10930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_10_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_12_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_10_cordic_atan_w_valuenode_10_w_range10929w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_10_cordic_atan_w_valuenode_12_w_range10927w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop2 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_10_cordic_atan_w_lg_w_lg_indexbit10930w10931w(i) <= wire_cata_10_cordic_atan_w_lg_indexbit10930w(0) AND wire_cata_10_cordic_atan_w_valuenode_10_w_range10929w(i);
	END GENERATE loop2;
	loop3 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_10_cordic_atan_w_lg_indexbit10928w(i) <= indexbit AND wire_cata_10_cordic_atan_w_valuenode_12_w_range10927w(i);
	END GENERATE loop3;
	wire_cata_10_cordic_atan_w_lg_indexbit10930w(0) <= NOT indexbit;
	arctan <= (wire_cata_10_cordic_atan_w_lg_w_lg_indexbit10930w10931w OR wire_cata_10_cordic_atan_w_lg_indexbit10928w);
	valuenode_10_w <= "000000000000111111111111111111111010101010101011";
	valuenode_12_w <= "000000000000001111111111111111111111111010101011";
	wire_cata_10_cordic_atan_w_valuenode_10_w_range10929w <= valuenode_10_w(47 DOWNTO 14);
	wire_cata_10_cordic_atan_w_valuenode_12_w_range10927w <= valuenode_12_w(45 DOWNTO 12);

 END RTL; --mysincos_altfp_sincos_cordic_atan_h9b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" indexpoint=2 START=11 WIDTH=34 arctan indexbit
--VERSION_BEGIN 13.0 cbx_altfp_sincos 2013:06:12:18:03:43:SJ cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_clshift 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altfp_sincos_cordic_atan_i9b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END mysincos_altfp_sincos_cordic_atan_i9b;

 ARCHITECTURE RTL OF mysincos_altfp_sincos_cordic_atan_i9b IS

	 SIGNAL  wire_cata_11_cordic_atan_w_lg_w_lg_indexbit10936w10937w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_11_cordic_atan_w_lg_indexbit10934w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_11_cordic_atan_w_lg_indexbit10936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_11_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_13_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_11_cordic_atan_w_valuenode_11_w_range10935w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_11_cordic_atan_w_valuenode_13_w_range10933w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop4 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_11_cordic_atan_w_lg_w_lg_indexbit10936w10937w(i) <= wire_cata_11_cordic_atan_w_lg_indexbit10936w(0) AND wire_cata_11_cordic_atan_w_valuenode_11_w_range10935w(i);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_11_cordic_atan_w_lg_indexbit10934w(i) <= indexbit AND wire_cata_11_cordic_atan_w_valuenode_13_w_range10933w(i);
	END GENERATE loop5;
	wire_cata_11_cordic_atan_w_lg_indexbit10936w(0) <= NOT indexbit;
	arctan <= (wire_cata_11_cordic_atan_w_lg_w_lg_indexbit10936w10937w OR wire_cata_11_cordic_atan_w_lg_indexbit10934w);
	valuenode_11_w <= "000000000000011111111111111111111111010101010101";
	valuenode_13_w <= "000000000000000111111111111111111111111111010101";
	wire_cata_11_cordic_atan_w_valuenode_11_w_range10935w <= valuenode_11_w(47 DOWNTO 14);
	wire_cata_11_cordic_atan_w_valuenode_13_w_range10933w <= valuenode_13_w(45 DOWNTO 12);

 END RTL; --mysincos_altfp_sincos_cordic_atan_i9b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" indexpoint=2 START=12 WIDTH=34 arctan indexbit
--VERSION_BEGIN 13.0 cbx_altfp_sincos 2013:06:12:18:03:43:SJ cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_clshift 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altfp_sincos_cordic_atan_j9b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END mysincos_altfp_sincos_cordic_atan_j9b;

 ARCHITECTURE RTL OF mysincos_altfp_sincos_cordic_atan_j9b IS

	 SIGNAL  wire_cata_12_cordic_atan_w_lg_w_lg_indexbit10942w10943w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_12_cordic_atan_w_lg_indexbit10940w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_12_cordic_atan_w_lg_indexbit10942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_12_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_14_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_12_cordic_atan_w_valuenode_12_w_range10941w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_12_cordic_atan_w_valuenode_14_w_range10939w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop6 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_12_cordic_atan_w_lg_w_lg_indexbit10942w10943w(i) <= wire_cata_12_cordic_atan_w_lg_indexbit10942w(0) AND wire_cata_12_cordic_atan_w_valuenode_12_w_range10941w(i);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_12_cordic_atan_w_lg_indexbit10940w(i) <= indexbit AND wire_cata_12_cordic_atan_w_valuenode_14_w_range10939w(i);
	END GENERATE loop7;
	wire_cata_12_cordic_atan_w_lg_indexbit10942w(0) <= NOT indexbit;
	arctan <= (wire_cata_12_cordic_atan_w_lg_w_lg_indexbit10942w10943w OR wire_cata_12_cordic_atan_w_lg_indexbit10940w);
	valuenode_12_w <= "000000000000001111111111111111111111111010101011";
	valuenode_14_w <= "000000000000000011111111111111111111111111111011";
	wire_cata_12_cordic_atan_w_valuenode_12_w_range10941w <= valuenode_12_w(47 DOWNTO 14);
	wire_cata_12_cordic_atan_w_valuenode_14_w_range10939w <= valuenode_14_w(45 DOWNTO 12);

 END RTL; --mysincos_altfp_sincos_cordic_atan_j9b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" indexpoint=2 START=13 WIDTH=34 arctan indexbit
--VERSION_BEGIN 13.0 cbx_altfp_sincos 2013:06:12:18:03:43:SJ cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_clshift 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altfp_sincos_cordic_atan_k9b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END mysincos_altfp_sincos_cordic_atan_k9b;

 ARCHITECTURE RTL OF mysincos_altfp_sincos_cordic_atan_k9b IS

	 SIGNAL  wire_cata_13_cordic_atan_w_lg_w_lg_indexbit10948w10949w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_13_cordic_atan_w_lg_indexbit10946w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_13_cordic_atan_w_lg_indexbit10948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_13_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_15_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_13_cordic_atan_w_valuenode_13_w_range10947w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_13_cordic_atan_w_valuenode_15_w_range10945w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop8 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_13_cordic_atan_w_lg_w_lg_indexbit10948w10949w(i) <= wire_cata_13_cordic_atan_w_lg_indexbit10948w(0) AND wire_cata_13_cordic_atan_w_valuenode_13_w_range10947w(i);
	END GENERATE loop8;
	loop9 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_13_cordic_atan_w_lg_indexbit10946w(i) <= indexbit AND wire_cata_13_cordic_atan_w_valuenode_15_w_range10945w(i);
	END GENERATE loop9;
	wire_cata_13_cordic_atan_w_lg_indexbit10948w(0) <= NOT indexbit;
	arctan <= (wire_cata_13_cordic_atan_w_lg_w_lg_indexbit10948w10949w OR wire_cata_13_cordic_atan_w_lg_indexbit10946w);
	valuenode_13_w <= "000000000000000111111111111111111111111111010101";
	valuenode_15_w <= "000000000000000001111111111111111111111111111111";
	wire_cata_13_cordic_atan_w_valuenode_13_w_range10947w <= valuenode_13_w(47 DOWNTO 14);
	wire_cata_13_cordic_atan_w_valuenode_15_w_range10945w <= valuenode_15_w(45 DOWNTO 12);

 END RTL; --mysincos_altfp_sincos_cordic_atan_k9b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" indexpoint=2 START=1 WIDTH=34 arctan indexbit
--VERSION_BEGIN 13.0 cbx_altfp_sincos 2013:06:12:18:03:43:SJ cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_clshift 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altfp_sincos_cordic_atan_18b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END mysincos_altfp_sincos_cordic_atan_18b;

 ARCHITECTURE RTL OF mysincos_altfp_sincos_cordic_atan_18b IS

	 SIGNAL  wire_cata_1_cordic_atan_w_lg_w_lg_indexbit10954w10955w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_1_cordic_atan_w_lg_indexbit10952w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_1_cordic_atan_w_lg_indexbit10954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_1_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_3_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_1_cordic_atan_w_valuenode_1_w_range10953w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_1_cordic_atan_w_valuenode_3_w_range10951w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop10 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_1_cordic_atan_w_lg_w_lg_indexbit10954w10955w(i) <= wire_cata_1_cordic_atan_w_lg_indexbit10954w(0) AND wire_cata_1_cordic_atan_w_valuenode_1_w_range10953w(i);
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_1_cordic_atan_w_lg_indexbit10952w(i) <= indexbit AND wire_cata_1_cordic_atan_w_valuenode_3_w_range10951w(i);
	END GENERATE loop11;
	wire_cata_1_cordic_atan_w_lg_indexbit10954w(0) <= NOT indexbit;
	arctan <= (wire_cata_1_cordic_atan_w_lg_w_lg_indexbit10954w10955w OR wire_cata_1_cordic_atan_w_lg_indexbit10952w);
	valuenode_1_w <= "000111011010110001100111000001010110000110111011";
	valuenode_3_w <= "000001111111010101101110101001101010101100001100";
	wire_cata_1_cordic_atan_w_valuenode_1_w_range10953w <= valuenode_1_w(47 DOWNTO 14);
	wire_cata_1_cordic_atan_w_valuenode_3_w_range10951w <= valuenode_3_w(45 DOWNTO 12);

 END RTL; --mysincos_altfp_sincos_cordic_atan_18b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" indexpoint=2 START=2 WIDTH=34 arctan indexbit
--VERSION_BEGIN 13.0 cbx_altfp_sincos 2013:06:12:18:03:43:SJ cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_clshift 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altfp_sincos_cordic_atan_28b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END mysincos_altfp_sincos_cordic_atan_28b;

 ARCHITECTURE RTL OF mysincos_altfp_sincos_cordic_atan_28b IS

	 SIGNAL  wire_cata_2_cordic_atan_w_lg_w_lg_indexbit10960w10961w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_2_cordic_atan_w_lg_indexbit10958w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_2_cordic_atan_w_lg_indexbit10960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_2_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_4_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_2_cordic_atan_w_valuenode_2_w_range10959w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_2_cordic_atan_w_valuenode_4_w_range10957w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop12 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_2_cordic_atan_w_lg_w_lg_indexbit10960w10961w(i) <= wire_cata_2_cordic_atan_w_lg_indexbit10960w(0) AND wire_cata_2_cordic_atan_w_valuenode_2_w_range10959w(i);
	END GENERATE loop12;
	loop13 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_2_cordic_atan_w_lg_indexbit10958w(i) <= indexbit AND wire_cata_2_cordic_atan_w_valuenode_4_w_range10957w(i);
	END GENERATE loop13;
	wire_cata_2_cordic_atan_w_lg_indexbit10960w(0) <= NOT indexbit;
	arctan <= (wire_cata_2_cordic_atan_w_lg_w_lg_indexbit10960w10961w OR wire_cata_2_cordic_atan_w_lg_indexbit10958w);
	valuenode_2_w <= "000011111010110110111010111111001001011001000000";
	valuenode_4_w <= "000000111111111010101011011101101110010110100000";
	wire_cata_2_cordic_atan_w_valuenode_2_w_range10959w <= valuenode_2_w(47 DOWNTO 14);
	wire_cata_2_cordic_atan_w_valuenode_4_w_range10957w <= valuenode_4_w(45 DOWNTO 12);

 END RTL; --mysincos_altfp_sincos_cordic_atan_28b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" indexpoint=2 START=3 WIDTH=34 arctan indexbit
--VERSION_BEGIN 13.0 cbx_altfp_sincos 2013:06:12:18:03:43:SJ cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_clshift 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altfp_sincos_cordic_atan_38b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END mysincos_altfp_sincos_cordic_atan_38b;

 ARCHITECTURE RTL OF mysincos_altfp_sincos_cordic_atan_38b IS

	 SIGNAL  wire_cata_3_cordic_atan_w_lg_w_lg_indexbit10966w10967w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_3_cordic_atan_w_lg_indexbit10964w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_3_cordic_atan_w_lg_indexbit10966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_3_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_5_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_3_cordic_atan_w_valuenode_3_w_range10965w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_3_cordic_atan_w_valuenode_5_w_range10963w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop14 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_3_cordic_atan_w_lg_w_lg_indexbit10966w10967w(i) <= wire_cata_3_cordic_atan_w_lg_indexbit10966w(0) AND wire_cata_3_cordic_atan_w_valuenode_3_w_range10965w(i);
	END GENERATE loop14;
	loop15 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_3_cordic_atan_w_lg_indexbit10964w(i) <= indexbit AND wire_cata_3_cordic_atan_w_valuenode_5_w_range10963w(i);
	END GENERATE loop15;
	wire_cata_3_cordic_atan_w_lg_indexbit10966w(0) <= NOT indexbit;
	arctan <= (wire_cata_3_cordic_atan_w_lg_w_lg_indexbit10966w10967w OR wire_cata_3_cordic_atan_w_lg_indexbit10964w);
	valuenode_3_w <= "000001111111010101101110101001101010101100001100";
	valuenode_5_w <= "000000011111111111010101010110111011101010010111";
	wire_cata_3_cordic_atan_w_valuenode_3_w_range10965w <= valuenode_3_w(47 DOWNTO 14);
	wire_cata_3_cordic_atan_w_valuenode_5_w_range10963w <= valuenode_5_w(45 DOWNTO 12);

 END RTL; --mysincos_altfp_sincos_cordic_atan_38b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" indexpoint=2 START=4 WIDTH=34 arctan indexbit
--VERSION_BEGIN 13.0 cbx_altfp_sincos 2013:06:12:18:03:43:SJ cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_clshift 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altfp_sincos_cordic_atan_48b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END mysincos_altfp_sincos_cordic_atan_48b;

 ARCHITECTURE RTL OF mysincos_altfp_sincos_cordic_atan_48b IS

	 SIGNAL  wire_cata_4_cordic_atan_w_lg_w_lg_indexbit10972w10973w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_4_cordic_atan_w_lg_indexbit10970w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_4_cordic_atan_w_lg_indexbit10972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_4_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_6_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_4_cordic_atan_w_valuenode_4_w_range10971w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_4_cordic_atan_w_valuenode_6_w_range10969w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop16 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_4_cordic_atan_w_lg_w_lg_indexbit10972w10973w(i) <= wire_cata_4_cordic_atan_w_lg_indexbit10972w(0) AND wire_cata_4_cordic_atan_w_valuenode_4_w_range10971w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_4_cordic_atan_w_lg_indexbit10970w(i) <= indexbit AND wire_cata_4_cordic_atan_w_valuenode_6_w_range10969w(i);
	END GENERATE loop17;
	wire_cata_4_cordic_atan_w_lg_indexbit10972w(0) <= NOT indexbit;
	arctan <= (wire_cata_4_cordic_atan_w_lg_w_lg_indexbit10972w10973w OR wire_cata_4_cordic_atan_w_lg_indexbit10970w);
	valuenode_4_w <= "000000111111111010101011011101101110010110100000";
	valuenode_6_w <= "000000001111111111111010101010101101110111011100";
	wire_cata_4_cordic_atan_w_valuenode_4_w_range10971w <= valuenode_4_w(47 DOWNTO 14);
	wire_cata_4_cordic_atan_w_valuenode_6_w_range10969w <= valuenode_6_w(45 DOWNTO 12);

 END RTL; --mysincos_altfp_sincos_cordic_atan_48b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" indexpoint=2 START=5 WIDTH=34 arctan indexbit
--VERSION_BEGIN 13.0 cbx_altfp_sincos 2013:06:12:18:03:43:SJ cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_clshift 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altfp_sincos_cordic_atan_58b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END mysincos_altfp_sincos_cordic_atan_58b;

 ARCHITECTURE RTL OF mysincos_altfp_sincos_cordic_atan_58b IS

	 SIGNAL  wire_cata_5_cordic_atan_w_lg_w_lg_indexbit10978w10979w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_5_cordic_atan_w_lg_indexbit10976w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_5_cordic_atan_w_lg_indexbit10978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_5_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_7_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_5_cordic_atan_w_valuenode_5_w_range10977w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_5_cordic_atan_w_valuenode_7_w_range10975w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop18 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_5_cordic_atan_w_lg_w_lg_indexbit10978w10979w(i) <= wire_cata_5_cordic_atan_w_lg_indexbit10978w(0) AND wire_cata_5_cordic_atan_w_valuenode_5_w_range10977w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_5_cordic_atan_w_lg_indexbit10976w(i) <= indexbit AND wire_cata_5_cordic_atan_w_valuenode_7_w_range10975w(i);
	END GENERATE loop19;
	wire_cata_5_cordic_atan_w_lg_indexbit10978w(0) <= NOT indexbit;
	arctan <= (wire_cata_5_cordic_atan_w_lg_w_lg_indexbit10978w10979w OR wire_cata_5_cordic_atan_w_lg_indexbit10976w);
	valuenode_5_w <= "000000011111111111010101010110111011101010010111";
	valuenode_7_w <= "000000000111111111111111010101010101011011101111";
	wire_cata_5_cordic_atan_w_valuenode_5_w_range10977w <= valuenode_5_w(47 DOWNTO 14);
	wire_cata_5_cordic_atan_w_valuenode_7_w_range10975w <= valuenode_7_w(45 DOWNTO 12);

 END RTL; --mysincos_altfp_sincos_cordic_atan_58b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" indexpoint=2 START=6 WIDTH=34 arctan indexbit
--VERSION_BEGIN 13.0 cbx_altfp_sincos 2013:06:12:18:03:43:SJ cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_clshift 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altfp_sincos_cordic_atan_68b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END mysincos_altfp_sincos_cordic_atan_68b;

 ARCHITECTURE RTL OF mysincos_altfp_sincos_cordic_atan_68b IS

	 SIGNAL  wire_cata_6_cordic_atan_w_lg_w_lg_indexbit10984w10985w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_6_cordic_atan_w_lg_indexbit10982w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_6_cordic_atan_w_lg_indexbit10984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_6_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_8_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_6_cordic_atan_w_valuenode_6_w_range10983w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_6_cordic_atan_w_valuenode_8_w_range10981w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop20 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_6_cordic_atan_w_lg_w_lg_indexbit10984w10985w(i) <= wire_cata_6_cordic_atan_w_lg_indexbit10984w(0) AND wire_cata_6_cordic_atan_w_valuenode_6_w_range10983w(i);
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_6_cordic_atan_w_lg_indexbit10982w(i) <= indexbit AND wire_cata_6_cordic_atan_w_valuenode_8_w_range10981w(i);
	END GENERATE loop21;
	wire_cata_6_cordic_atan_w_lg_indexbit10984w(0) <= NOT indexbit;
	arctan <= (wire_cata_6_cordic_atan_w_lg_w_lg_indexbit10984w10985w OR wire_cata_6_cordic_atan_w_lg_indexbit10982w);
	valuenode_6_w <= "000000001111111111111010101010101101110111011100";
	valuenode_8_w <= "000000000011111111111111111010101010101010110111";
	wire_cata_6_cordic_atan_w_valuenode_6_w_range10983w <= valuenode_6_w(47 DOWNTO 14);
	wire_cata_6_cordic_atan_w_valuenode_8_w_range10981w <= valuenode_8_w(45 DOWNTO 12);

 END RTL; --mysincos_altfp_sincos_cordic_atan_68b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" indexpoint=2 START=7 WIDTH=34 arctan indexbit
--VERSION_BEGIN 13.0 cbx_altfp_sincos 2013:06:12:18:03:43:SJ cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_clshift 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altfp_sincos_cordic_atan_78b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END mysincos_altfp_sincos_cordic_atan_78b;

 ARCHITECTURE RTL OF mysincos_altfp_sincos_cordic_atan_78b IS

	 SIGNAL  wire_cata_7_cordic_atan_w_lg_w_lg_indexbit10990w10991w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_7_cordic_atan_w_lg_indexbit10988w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_7_cordic_atan_w_lg_indexbit10990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_7_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_9_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_7_cordic_atan_w_valuenode_7_w_range10989w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_7_cordic_atan_w_valuenode_9_w_range10987w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop22 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_7_cordic_atan_w_lg_w_lg_indexbit10990w10991w(i) <= wire_cata_7_cordic_atan_w_lg_indexbit10990w(0) AND wire_cata_7_cordic_atan_w_valuenode_7_w_range10989w(i);
	END GENERATE loop22;
	loop23 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_7_cordic_atan_w_lg_indexbit10988w(i) <= indexbit AND wire_cata_7_cordic_atan_w_valuenode_9_w_range10987w(i);
	END GENERATE loop23;
	wire_cata_7_cordic_atan_w_lg_indexbit10990w(0) <= NOT indexbit;
	arctan <= (wire_cata_7_cordic_atan_w_lg_w_lg_indexbit10990w10991w OR wire_cata_7_cordic_atan_w_lg_indexbit10988w);
	valuenode_7_w <= "000000000111111111111111010101010101011011101111";
	valuenode_9_w <= "000000000001111111111111111111010101010101010110";
	wire_cata_7_cordic_atan_w_valuenode_7_w_range10989w <= valuenode_7_w(47 DOWNTO 14);
	wire_cata_7_cordic_atan_w_valuenode_9_w_range10987w <= valuenode_9_w(45 DOWNTO 12);

 END RTL; --mysincos_altfp_sincos_cordic_atan_78b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" indexpoint=2 START=8 WIDTH=34 arctan indexbit
--VERSION_BEGIN 13.0 cbx_altfp_sincos 2013:06:12:18:03:43:SJ cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_clshift 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altfp_sincos_cordic_atan_88b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END mysincos_altfp_sincos_cordic_atan_88b;

 ARCHITECTURE RTL OF mysincos_altfp_sincos_cordic_atan_88b IS

	 SIGNAL  wire_cata_8_cordic_atan_w_lg_w_lg_indexbit10996w10997w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_8_cordic_atan_w_lg_indexbit10994w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_8_cordic_atan_w_lg_indexbit10996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_10_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_8_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_8_cordic_atan_w_valuenode_10_w_range10993w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_8_cordic_atan_w_valuenode_8_w_range10995w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop24 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_8_cordic_atan_w_lg_w_lg_indexbit10996w10997w(i) <= wire_cata_8_cordic_atan_w_lg_indexbit10996w(0) AND wire_cata_8_cordic_atan_w_valuenode_8_w_range10995w(i);
	END GENERATE loop24;
	loop25 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_8_cordic_atan_w_lg_indexbit10994w(i) <= indexbit AND wire_cata_8_cordic_atan_w_valuenode_10_w_range10993w(i);
	END GENERATE loop25;
	wire_cata_8_cordic_atan_w_lg_indexbit10996w(0) <= NOT indexbit;
	arctan <= (wire_cata_8_cordic_atan_w_lg_w_lg_indexbit10996w10997w OR wire_cata_8_cordic_atan_w_lg_indexbit10994w);
	valuenode_10_w <= "000000000000111111111111111111111010101010101011";
	valuenode_8_w <= "000000000011111111111111111010101010101010110111";
	wire_cata_8_cordic_atan_w_valuenode_10_w_range10993w <= valuenode_10_w(45 DOWNTO 12);
	wire_cata_8_cordic_atan_w_valuenode_8_w_range10995w <= valuenode_8_w(47 DOWNTO 14);

 END RTL; --mysincos_altfp_sincos_cordic_atan_88b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" indexpoint=2 START=9 WIDTH=34 arctan indexbit
--VERSION_BEGIN 13.0 cbx_altfp_sincos 2013:06:12:18:03:43:SJ cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_clshift 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altfp_sincos_cordic_atan_98b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END mysincos_altfp_sincos_cordic_atan_98b;

 ARCHITECTURE RTL OF mysincos_altfp_sincos_cordic_atan_98b IS

	 SIGNAL  wire_cata_9_cordic_atan_w_lg_w_lg_indexbit11002w11003w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_9_cordic_atan_w_lg_indexbit11000w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_9_cordic_atan_w_lg_indexbit11002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_11_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_9_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_9_cordic_atan_w_valuenode_11_w_range10999w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_9_cordic_atan_w_valuenode_9_w_range11001w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop26 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_9_cordic_atan_w_lg_w_lg_indexbit11002w11003w(i) <= wire_cata_9_cordic_atan_w_lg_indexbit11002w(0) AND wire_cata_9_cordic_atan_w_valuenode_9_w_range11001w(i);
	END GENERATE loop26;
	loop27 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_9_cordic_atan_w_lg_indexbit11000w(i) <= indexbit AND wire_cata_9_cordic_atan_w_valuenode_11_w_range10999w(i);
	END GENERATE loop27;
	wire_cata_9_cordic_atan_w_lg_indexbit11002w(0) <= NOT indexbit;
	arctan <= (wire_cata_9_cordic_atan_w_lg_w_lg_indexbit11002w11003w OR wire_cata_9_cordic_atan_w_lg_indexbit11000w);
	valuenode_11_w <= "000000000000011111111111111111111111010101010101";
	valuenode_9_w <= "000000000001111111111111111111010101010101010110";
	wire_cata_9_cordic_atan_w_valuenode_11_w_range10999w <= valuenode_11_w(45 DOWNTO 12);
	wire_cata_9_cordic_atan_w_valuenode_9_w_range11001w <= valuenode_9_w(47 DOWNTO 14);

 END RTL; --mysincos_altfp_sincos_cordic_atan_98b


--altfp_sincos_cordic_start CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" WIDTH=34 index value
--VERSION_BEGIN 13.0 cbx_altfp_sincos 2013:06:12:18:03:43:SJ cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_clshift 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.lpm_components.all;

--synthesis_resources = lpm_mux 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altfp_sincos_cordic_start_339 IS 
	 PORT 
	 ( 
		 index	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => '0');
		 value	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0)
	 ); 
 END mysincos_altfp_sincos_cordic_start_339;

 ARCHITECTURE RTL OF mysincos_altfp_sincos_cordic_start_339 IS

	 SIGNAL  wire_mux1_data	:	STD_LOGIC_VECTOR (543 DOWNTO 0);
	 SIGNAL  wire_mux1_data_2d	:	STD_LOGIC_2D(15 DOWNTO 0, 33 DOWNTO 0);
	 SIGNAL  wire_mux1_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  valuenode_0_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_10_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_11_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_12_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_13_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_14_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_15_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_1_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_2_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_3_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_4_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_5_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_6_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_7_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_8_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_9_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
 BEGIN

	value <= wire_mux1_result;
	valuenode_0_w <= "001001101101110100111011011010100001";
	valuenode_10_w <= "001111111111111111111101010101010101";
	valuenode_11_w <= "001111111111111111111111010101010101";
	valuenode_12_w <= "001111111111111111111111111101010101";
	valuenode_13_w <= "001111111111111111111111110101010101";
	valuenode_14_w <= "001111111111111111111111111111110101";
	valuenode_15_w <= "001111111111111111111111111111010101";
	valuenode_1_w <= "001101101111011001010110110001011010";
	valuenode_2_w <= "001111010111001100011101111111111011";
	valuenode_3_w <= "001111110101011101000011101100100100";
	valuenode_4_w <= "001111111101010101110100100001100000";
	valuenode_5_w <= "001111111111010101010111010010011001";
	valuenode_6_w <= "001111111111110101010101011101001010";
	valuenode_7_w <= "001111111111111101010101010101110101";
	valuenode_8_w <= "001111111111111111010101010101010111";
	valuenode_9_w <= "001111111111111111110101010101010101";
	wire_mux1_data <= ( valuenode_15_w(35 DOWNTO 2) & valuenode_14_w(35 DOWNTO 2) & valuenode_13_w(35 DOWNTO 2) & valuenode_12_w(35 DOWNTO 2) & valuenode_11_w(35 DOWNTO 2) & valuenode_10_w(35 DOWNTO 2) & valuenode_9_w(35 DOWNTO 2) & valuenode_8_w(35 DOWNTO 2) & valuenode_7_w(35 DOWNTO 2) & valuenode_6_w(35 DOWNTO 2) & valuenode_5_w(35 DOWNTO 2) & valuenode_4_w(35 DOWNTO 2) & valuenode_3_w(35 DOWNTO 2) & valuenode_2_w(35 DOWNTO 2) & valuenode_1_w(35 DOWNTO 2) & valuenode_0_w(35 DOWNTO 2));
	loop28 : FOR i IN 0 TO 15 GENERATE
		loop29 : FOR j IN 0 TO 33 GENERATE
			wire_mux1_data_2d(i, j) <= wire_mux1_data(i*34+j);
		END GENERATE loop29;
	END GENERATE loop28;
	mux1 :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 16,
		LPM_WIDTH => 34,
		LPM_WIDTHS => 4
	  )
	  PORT MAP ( 
		data => wire_mux1_data_2d,
		result => wire_mux1_result,
		sel => index
	  );

 END RTL; --mysincos_altfp_sincos_cordic_start_339

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 39 lpm_mult 1 lpm_mux 1 reg 1598 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altfp_sincos_cordic_m_a8e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 indexbit	:	IN  STD_LOGIC := '0';
		 radians	:	IN  STD_LOGIC_VECTOR (33 DOWNTO 0) := (OTHERS => '0');
		 sincos	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 sincosbit	:	IN  STD_LOGIC := '0'
	 ); 
 END mysincos_altfp_sincos_cordic_m_a8e;

 ARCHITECTURE RTL OF mysincos_altfp_sincos_cordic_m_a8e IS

	 SIGNAL  wire_cata_0_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_10_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_11_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_12_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_13_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_1_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_2_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_3_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_4_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_5_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_6_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_7_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_8_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_9_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cxs_value	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL	 cdaff_0	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cdaff_1	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cdaff_2	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 indexbitff	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_indexbitff_w_lg_w_q_range581w681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range610w8591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range613w9393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range616w10190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range10749w10754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range583w1148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range586w1995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range589w2837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range592w3674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range595w4506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range598w5333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range601w6155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range604w6972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range607w7784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range10749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 sincosbitff	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_sincosbitff_w_lg_w_q_range668w10739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_sincosbitff_w_lg_w_q_range10746w10747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_sincosbitff_w_q_range668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_sincosbitff_w_q_range10746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 sincosff	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_0	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range678w682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range721w734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range721w723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range726w739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range726w728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range731w744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range731w733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range736w749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range736w738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range741w754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range741w743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range746w759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range746w748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range751w764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range751w753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range756w769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range756w758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range761w774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range761w763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range766w779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range766w768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range686w689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range771w784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range771w773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range776w789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range776w778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range781w794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range781w783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range786w799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range786w788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range791w804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range791w793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range796w809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range796w798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range801w814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range801w803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range806w819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range806w808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range811w824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range811w813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range816w829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range816w818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range677w694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range677w680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range821w834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range821w823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range826w839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range826w828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range831w842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range831w833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range836w838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range685w699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range685w688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range691w704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range691w693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range696w709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range696w698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range701w714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range701w703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range706w719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range706w708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range711w724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range711w713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range716w729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range716w718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range836w844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range678w682w683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range721w734w735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range726w739w740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range731w744w745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range736w749w750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range741w754w755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range746w759w760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range751w764w765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range756w769w770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range761w774w775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range766w779w780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range686w689w690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range771w784w785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range776w789w790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range781w794w795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range786w799w800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range791w804w805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range796w809w810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range801w814w815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range806w819w820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range811w824w825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range816w829w830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range677w694w695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range821w834w835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range826w839w840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range685w699w700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range691w704w705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range696w709w710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range701w714w715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range706w719w720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range711w724w725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range716w729w730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 x_pipeff_1	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_10	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_11	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_12	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_13	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_x_pipeff_13_w_lg_q10744w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_13_w_lg_q10741w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL	 x_pipeff_2	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_3	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_4	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_5	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_6	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_7	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_8	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_9	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 y_pipeff_0	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 y_pipeff_1	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range913w915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range919w921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range925w927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range931w933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range937w939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range943w945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range949w951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range955w957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range961w963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range967w969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range860w862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range973w975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range979w981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range985w987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range991w993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range997w999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range1003w1005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range1009w1011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range1015w1017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range1021w1023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range1027w1029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range865w867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range1033w1035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range1039w1041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range1045w1047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range845w847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range871w873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range877w879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range883w885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range889w891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range895w897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range901w903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range907w909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range1003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range1009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range1015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range1021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range1027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range1033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range1039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range1045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_10	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8384w8386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8389w8391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8395w8397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8401w8403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8407w8409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8413w8415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8419w8421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8425w8427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8431w8433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8437w8439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8443w8445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8449w8451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8455w8457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8461w8463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8467w8469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8473w8475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8479w8481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8485w8487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8491w8493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8497w8499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8503w8505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8509w8511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8515w8517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8333w8335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_11	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9195w9197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9200w9202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9206w9208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9212w9214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9218w9220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9224w9226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9230w9232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9236w9238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9242w9244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9248w9250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9254w9256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9260w9262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9266w9268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9272w9274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9278w9280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9284w9286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9290w9292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9296w9298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9302w9304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9308w9310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9314w9316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9320w9322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9140w9142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_12	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10001w10003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10006w10008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10012w10014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10018w10020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10024w10026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10030w10032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10036w10038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10042w10044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10048w10050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10054w10056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10060w10062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10066w10068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10072w10074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10078w10080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10084w10086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10090w10092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10096w10098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10102w10104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10108w10110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10114w10116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10120w10122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range9942w9944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range9942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_13	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_13_w_lg_q10740w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_13_w_lg_q10743w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL	 y_pipeff_2	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1763w1765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1769w1771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1775w1777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1781w1783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1787w1789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1793w1795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1799w1801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1805w1807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1811w1813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1817w1819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1823w1825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1829w1831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1835w1837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1841w1843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1847w1849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1853w1855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1859w1861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1865w1867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1871w1873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1877w1879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1716w1718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1883w1885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1889w1891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1895w1897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1697w1699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1721w1723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1727w1729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1733w1735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1739w1741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1745w1747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1751w1753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1757w1759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_3	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2608w2610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2614w2616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2620w2622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2626w2628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2632w2634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2638w2640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2644w2646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2650w2652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2656w2658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2662w2664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2668w2670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2674w2676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2680w2682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2686w2688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2692w2694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2698w2700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2704w2706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2710w2712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2716w2718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2722w2724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2728w2730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2734w2736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2740w2742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2544w2546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2567w2569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2572w2574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2578w2580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2584w2586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2590w2592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2596w2598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2602w2604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_4	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3448w3450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3454w3456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3460w3462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3466w3468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3472w3474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3478w3480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3484w3486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3490w3492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3496w3498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3502w3504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3508w3510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3514w3516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3520w3522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3526w3528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3532w3534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3538w3540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3544w3546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3550w3552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3556w3558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3562w3564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3568w3570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3574w3576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3580w3582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3386w3388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3413w3415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3418w3420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3424w3426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3430w3432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3436w3438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3442w3444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_5	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4283w4285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4289w4291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4295w4297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4301w4303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4307w4309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4313w4315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4319w4321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4325w4327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4331w4333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4337w4339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4343w4345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4349w4351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4355w4357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4361w4363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4367w4369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4373w4375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4379w4381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4385w4387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4391w4393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4397w4399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4403w4405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4409w4411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4415w4417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4223w4225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4254w4256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4259w4261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4265w4267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4271w4273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4277w4279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_6	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5113w5115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5119w5121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5125w5127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5131w5133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5137w5139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5143w5145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5149w5151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5155w5157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5161w5163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5167w5169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5173w5175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5179w5181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5185w5187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5191w5193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5197w5199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5203w5205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5209w5211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5215w5217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5221w5223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5227w5229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5233w5235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5239w5241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5245w5247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5055w5057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5090w5092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5095w5097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5101w5103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5107w5109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_7	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5938w5940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5944w5946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5950w5952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5956w5958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5962w5964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5968w5970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5974w5976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5980w5982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5986w5988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5992w5994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5998w6000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6004w6006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6010w6012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6016w6018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6022w6024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6028w6030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6034w6036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6040w6042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6046w6048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6052w6054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6058w6060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6064w6066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6070w6072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5882w5884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5921w5923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5926w5928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5932w5934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_8	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6758w6760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6764w6766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6770w6772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6776w6778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6782w6784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6788w6790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6794w6796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6800w6802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6806w6808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6812w6814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6818w6820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6824w6826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6830w6832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6836w6838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6842w6844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6848w6850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6854w6856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6860w6862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6866w6868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6872w6874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6878w6880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6884w6886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6890w6892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6704w6706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6747w6749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6752w6754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_9	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7573w7575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7579w7581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7585w7587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7591w7593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7597w7599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7603w7605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7609w7611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7615w7617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7621w7623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7627w7629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7633w7635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7639w7641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7645w7647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7651w7653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7657w7659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7663w7665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7669w7671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7675w7677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7681w7683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7687w7689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7693w7695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7699w7701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7705w7707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7521w7523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7568w7570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_0	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 z_pipeff_1	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_1_w_q_range1421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_10	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_10_w_q_range8864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_11	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_11_w_q_range9666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_12	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_12_w_q_range10463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_13	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 z_pipeff_2	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_2_w_q_range2268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_3	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_3_w_q_range3110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_4	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_4_w_q_range3947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_5	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_5_w_q_range4779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_6	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_6_w_q_range5606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_7	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_7_w_q_range6428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_8	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_8_w_q_range7245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_9	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_9_w_q_range8057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_sincos_add_cin	:	STD_LOGIC;
	 SIGNAL  wire_sincos_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_10_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_11_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_12_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_13_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_2_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_3_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_4_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_5_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_6_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_7_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_8_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_9_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipeff1_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_10_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_11_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_12_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_13_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_2_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_3_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_4_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_5_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_6_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_7_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_8_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_9_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipeff1_sub_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_10_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_11_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_12_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_13_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_2_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_3_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_4_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_5_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_6_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_7_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_8_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_9_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cmx_result	:	STD_LOGIC_VECTOR (67 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_indexpointnum_w409w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10751w10755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10794w10807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10794w10796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10799w10812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10799w10801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10804w10817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10804w10806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10809w10822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10809w10811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10814w10827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10814w10816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10819w10832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10819w10821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10824w10837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10824w10826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10829w10842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10829w10831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10834w10847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10834w10836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10839w10852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10839w10841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10759w10762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10844w10857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10844w10846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10849w10862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10849w10851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10854w10867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10854w10856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10859w10872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10859w10861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10864w10877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10864w10866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10869w10882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10869w10871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10874w10887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10874w10876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10879w10892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10879w10881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10884w10897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10884w10886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10889w10902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10889w10891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10750w10767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10750w10753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10894w10907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10894w10896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10899w10912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10899w10901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10904w10915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10904w10906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10909w10918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10909w10911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10758w10772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10758w10761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10764w10777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10764w10766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10769w10782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10769w10771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10774w10787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10774w10776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10779w10792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10779w10781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10784w10797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10784w10786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10789w10802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10789w10791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range410w413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range410w420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range458w461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range458w470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range463w466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range463w475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range468w471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range468w480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range473w476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range473w485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range478w481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range478w490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range483w486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range483w495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range488w491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range488w500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range493w496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range493w505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range498w501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range498w510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range503w506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range503w515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range415w417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range415w425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range508w511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range508w520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range513w516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range513w525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range518w521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range518w530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range523w526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range523w535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range528w531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range528w540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range533w536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range533w545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range538w541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range538w550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range543w546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range543w555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range548w551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range548w560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range553w556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range553w565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range418w421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range418w430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range558w561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range558w570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range563w566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range563w575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range568w571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range573w576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range423w426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range423w435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range428w431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range428w440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range433w436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range433w445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range438w441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range438w450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range443w446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range443w455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range448w451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range448w460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range453w456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range453w465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7569w7785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7628w7867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7634w7875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7640w7883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7646w7891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7652w7899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7658w7907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7664w7915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7670w7923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7676w7931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7682w7939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7574w7795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7688w7947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7694w7955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7700w7963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7706w7971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7711w7979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7522w7987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7528w7995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7530w8003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7532w8011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7534w8019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7580w7803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7536w8027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7538w8035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7540w8043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7542w8051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7586w7811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7592w7819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7598w7827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7604w7835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7610w7843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7616w7851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7622w7859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8385w8592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8444w8674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8450w8682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8456w8690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8462w8698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8468w8706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8474w8714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8480w8722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8486w8730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8492w8738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8498w8746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8390w8602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8504w8754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8510w8762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8516w8770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8521w8778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8334w8786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8340w8794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8342w8802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8344w8810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8346w8818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8348w8826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8396w8610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8350w8834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8352w8842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8354w8850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8356w8858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8402w8618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8408w8626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8414w8634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8420w8642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8426w8650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8432w8658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8438w8666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9196w9394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9255w9476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9261w9484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9267w9492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9273w9500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9279w9508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9285w9516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9291w9524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9297w9532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9303w9540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9309w9548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9201w9404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9315w9556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9321w9564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9326w9572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9141w9580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9147w9588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9149w9596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9151w9604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9153w9612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9155w9620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9157w9628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9207w9412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9159w9636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9161w9644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9163w9652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9165w9660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9213w9420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9219w9428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9225w9436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9231w9444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9237w9452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9243w9460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9249w9468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10002w10191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10061w10273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10067w10281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10073w10289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10079w10297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10085w10305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10091w10313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10097w10321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10103w10329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10109w10337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10115w10345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10007w10201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10121w10353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10126w10361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9943w10369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9949w10377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9951w10385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9953w10393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9955w10401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9957w10409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9959w10417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9961w10425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10013w10209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9963w10433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9965w10441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9967w10449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9969w10457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10019w10217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10025w10225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10031w10233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10037w10241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10043w10249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10049w10257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10055w10265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range861w1149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range920w1231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range926w1239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range932w1247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range938w1255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range944w1263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range950w1271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range956w1279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range962w1287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range968w1295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range974w1303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range866w1159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range980w1311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range986w1319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range992w1327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range998w1335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1004w1343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1010w1351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1016w1359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1022w1367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1028w1375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1034w1383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range872w1167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1040w1391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1046w1399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1051w1407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range846w1415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range878w1175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range884w1183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range890w1191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range896w1199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range902w1207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range908w1215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range914w1223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1717w1996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1776w2078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1782w2086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1788w2094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1794w2102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1800w2110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1806w2118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1812w2126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1818w2134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1824w2142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1830w2150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1722w2006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1836w2158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1842w2166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1848w2174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1854w2182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1860w2190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1866w2198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1872w2206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1878w2214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1884w2222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1890w2230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1728w2014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1896w2238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1901w2246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1698w2254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1704w2262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1734w2022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1740w2030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1746w2038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1752w2046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1758w2054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1764w2062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1770w2070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2568w2838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2627w2920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2633w2928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2639w2936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2645w2944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2651w2952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2657w2960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2663w2968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2669w2976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2675w2984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2681w2992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2573w2848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2687w3000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2693w3008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2699w3016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2705w3024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2711w3032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2717w3040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2723w3048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2729w3056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2735w3064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2741w3072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2579w2856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2746w3080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2545w3088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2551w3096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2553w3104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2585w2864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2591w2872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2597w2880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2603w2888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2609w2896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2615w2904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2621w2912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3414w3675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3473w3757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3479w3765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3485w3773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3491w3781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3497w3789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3503w3797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3509w3805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3515w3813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3521w3821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3527w3829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3419w3685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3533w3837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3539w3845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3545w3853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3551w3861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3557w3869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3563w3877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3569w3885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3575w3893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3581w3901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3586w3909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3425w3693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3387w3917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3393w3925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3395w3933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3397w3941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3431w3701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3437w3709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3443w3717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3449w3725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3455w3733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3461w3741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3467w3749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4255w4507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4314w4589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4320w4597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4326w4605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4332w4613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4338w4621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4344w4629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4350w4637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4356w4645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4362w4653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4368w4661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4260w4517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4374w4669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4380w4677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4386w4685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4392w4693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4398w4701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4404w4709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4410w4717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4416w4725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4421w4733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4224w4741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4266w4525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4230w4749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4232w4757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4234w4765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4236w4773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4272w4533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4278w4541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4284w4549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4290w4557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4296w4565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4302w4573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4308w4581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5091w5334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5150w5416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5156w5424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5162w5432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5168w5440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5174w5448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5180w5456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5186w5464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5192w5472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5198w5480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5204w5488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5096w5344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5210w5496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5216w5504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5222w5512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5228w5520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5234w5528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5240w5536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5246w5544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5251w5552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5056w5560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5062w5568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5102w5352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5064w5576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5066w5584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5068w5592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5070w5600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5108w5360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5114w5368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5120w5376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5126w5384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5132w5392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5138w5400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5144w5408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5922w6156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5981w6238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5987w6246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5993w6254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5999w6262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6005w6270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6011w6278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6017w6286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6023w6294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6029w6302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6035w6310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5927w6166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6041w6318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6047w6326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6053w6334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6059w6342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6065w6350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6071w6358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6076w6366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5883w6374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5889w6382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5891w6390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5933w6174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5893w6398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5895w6406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5897w6414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5899w6422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5939w6182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5945w6190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5951w6198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5957w6206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5963w6214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5969w6222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5975w6230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6748w6973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6807w7055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6813w7063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6819w7071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6825w7079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6831w7087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6837w7095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6843w7103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6849w7111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6855w7119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6861w7127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6753w6983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6867w7135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6873w7143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6879w7151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6885w7159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6891w7167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6896w7175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6705w7183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6711w7191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6713w7199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6715w7207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6759w6991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6717w7215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6719w7223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6721w7231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6723w7239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6765w6999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6771w7007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6777w7015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6783w7023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6789w7031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6795w7039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6801w7047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7714w7783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7743w7866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7746w7874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7749w7882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7752w7890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7755w7898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7758w7906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7761w7914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7764w7922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7767w7930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7770w7938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7716w7794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7773w7946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7776w7954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7779w7962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7544w7970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7548w7978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7550w7986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7552w7994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7554w8002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7556w8010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7558w8018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7719w7802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7560w8026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7562w8034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7564w8042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7566w8050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7722w7810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7725w7818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7728w7826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7731w7834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7734w7842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7737w7850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7740w7858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8524w8590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8553w8673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8556w8681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8559w8689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8562w8697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8565w8705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8568w8713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8571w8721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8574w8729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8577w8737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8580w8745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8526w8601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8583w8753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8586w8761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8358w8769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8362w8777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8364w8785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8366w8793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8368w8801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8370w8809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8372w8817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8374w8825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8529w8609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8376w8833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8378w8841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8380w8849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8382w8857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8532w8617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8535w8625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8538w8633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8541w8641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8544w8649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8547w8657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8550w8665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9329w9392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9358w9475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9361w9483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9364w9491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9367w9499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9370w9507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9373w9515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9376w9523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9379w9531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9382w9539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9385w9547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9331w9403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9388w9555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9167w9563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9171w9571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9173w9579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9175w9587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9177w9595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9179w9603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9181w9611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9183w9619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9185w9627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9334w9411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9187w9635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9189w9643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9191w9651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9193w9659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9337w9419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9340w9427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9343w9435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9346w9443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9349w9451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9352w9459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9355w9467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10129w10189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10158w10272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10161w10280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10164w10288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10167w10296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10170w10304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10173w10312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10176w10320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10179w10328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10182w10336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10185w10344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10131w10200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9971w10352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9975w10360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9977w10368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9979w10376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9981w10384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9983w10392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9985w10400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9987w10408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9989w10416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9991w10424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10134w10208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9993w10432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9995w10440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9997w10448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9999w10456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10137w10216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10140w10224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10143w10232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10146w10240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10149w10248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10152w10256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10155w10264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1054w1147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1083w1230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1086w1238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1089w1246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1092w1254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1095w1262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1098w1270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1101w1278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1104w1286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1107w1294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1110w1302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1056w1158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1113w1310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1116w1318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1119w1326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1122w1334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1125w1342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1128w1350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1131w1358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1134w1366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1137w1374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1140w1382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1059w1166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1143w1390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range852w1398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range856w1406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range858w1414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1062w1174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1065w1182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1068w1190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1071w1198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1074w1206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1077w1214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1080w1222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1904w1994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1933w2077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1936w2085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1939w2093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1942w2101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1945w2109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1948w2117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1951w2125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1954w2133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1957w2141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1960w2149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1906w2005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1963w2157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1966w2165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1969w2173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1972w2181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1975w2189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1978w2197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1981w2205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1984w2213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1987w2221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1990w2229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1909w2013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1706w2237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1710w2245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1712w2253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1714w2261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1912w2021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1915w2029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1918w2037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1921w2045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1924w2053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1927w2061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1930w2069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2749w2836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2778w2919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2781w2927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2784w2935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2787w2943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2790w2951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2793w2959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2796w2967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2799w2975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2802w2983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2805w2991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2751w2847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2808w2999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2811w3007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2814w3015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2817w3023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2820w3031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2823w3039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2826w3047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2829w3055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2832w3063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2555w3071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2754w2855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2559w3079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2561w3087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2563w3095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2565w3103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2757w2863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2760w2871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2763w2879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2766w2887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2769w2895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2772w2903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2775w2911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3589w3673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3618w3756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3621w3764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3624w3772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3627w3780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3630w3788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3633w3796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3636w3804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3639w3812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3642w3820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3645w3828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3591w3684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3648w3836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3651w3844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3654w3852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3657w3860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3660w3868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3663w3876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3666w3884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3669w3892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3399w3900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3403w3908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3594w3692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3405w3916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3407w3924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3409w3932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3411w3940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3597w3700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3600w3708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3603w3716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3606w3724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3609w3732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3612w3740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3615w3748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4424w4505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4453w4588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4456w4596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4459w4604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4462w4612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4465w4620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4468w4628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4471w4636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4474w4644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4477w4652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4480w4660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4426w4516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4483w4668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4486w4676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4489w4684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4492w4692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4495w4700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4498w4708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4501w4716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4238w4724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4242w4732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4244w4740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4429w4524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4246w4748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4248w4756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4250w4764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4252w4772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4432w4532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4435w4540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4438w4548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4441w4556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4444w4564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4447w4572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4450w4580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5254w5332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5283w5415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5286w5423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5289w5431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5292w5439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5295w5447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5298w5455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5301w5463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5304w5471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5307w5479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5310w5487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5256w5343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5313w5495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5316w5503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5319w5511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5322w5519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5325w5527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5328w5535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5072w5543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5076w5551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5078w5559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5080w5567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5259w5351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5082w5575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5084w5583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5086w5591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5088w5599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5262w5359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5265w5367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5268w5375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5271w5383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5274w5391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5277w5399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5280w5407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6079w6154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6108w6237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6111w6245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6114w6253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6117w6261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6120w6269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6123w6277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6126w6285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6129w6293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6132w6301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6135w6309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6081w6165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6138w6317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6141w6325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6144w6333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6147w6341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6150w6349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5901w6357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5905w6365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5907w6373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5909w6381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5911w6389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6084w6173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5913w6397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5915w6405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5917w6413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5919w6421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6087w6181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6090w6189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6093w6197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6096w6205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6099w6213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6102w6221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6105w6229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6899w6971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6928w7054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6931w7062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6934w7070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6937w7078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6940w7086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6943w7094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6946w7102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6949w7110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6952w7118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6955w7126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6901w6982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6958w7134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6961w7142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6964w7150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6967w7158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6725w7166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6729w7174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6731w7182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6733w7190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6735w7198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6737w7206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6904w6990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6739w7214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6741w7222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6743w7230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6745w7238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6907w6998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6910w7006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6913w7014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6916w7022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6919w7030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6922w7038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6925w7046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7572w7790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7631w7871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7637w7879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7643w7887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7649w7895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7655w7903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7661w7911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7667w7919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7673w7927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7679w7935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7685w7943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7577w7799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7691w7951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7697w7959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7703w7967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7709w7975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7712w7983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7526w7991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7529w7999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7531w8007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7533w8015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7535w8023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7583w7807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7537w8031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7539w8039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7541w8047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7543w8055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7589w7815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7595w7823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7601w7831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7607w7839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7613w7847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7619w7855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7625w7863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8388w8597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8447w8678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8453w8686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8459w8694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8465w8702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8471w8710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8477w8718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8483w8726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8489w8734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8495w8742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8501w8750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8393w8606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8507w8758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8513w8766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8519w8774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8522w8782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8338w8790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8341w8798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8343w8806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8345w8814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8347w8822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8349w8830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8399w8614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8351w8838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8353w8846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8355w8854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8357w8862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8405w8622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8411w8630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8417w8638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8423w8646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8429w8654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8435w8662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8441w8670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9199w9399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9258w9480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9264w9488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9270w9496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9276w9504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9282w9512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9288w9520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9294w9528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9300w9536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9306w9544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9312w9552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9204w9408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9318w9560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9324w9568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9327w9576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9145w9584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9148w9592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9150w9600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9152w9608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9154w9616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9156w9624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9158w9632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9210w9416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9160w9640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9162w9648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9164w9656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9166w9664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9216w9424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9222w9432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9228w9440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9234w9448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9240w9456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9246w9464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9252w9472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10005w10196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10064w10277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10070w10285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10076w10293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10082w10301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10088w10309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10094w10317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10100w10325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10106w10333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10112w10341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10118w10349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10010w10205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10124w10357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10127w10365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9947w10373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9950w10381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9952w10389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9954w10397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9956w10405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9958w10413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9960w10421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9962w10429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10016w10213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9964w10437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9966w10445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9968w10453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9970w10461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10022w10221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10028w10229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10034w10237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10040w10245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10046w10253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10052w10261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10058w10269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range864w1154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range923w1235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range929w1243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range935w1251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range941w1259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range947w1267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range953w1275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range959w1283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range965w1291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range971w1299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range977w1307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range869w1163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range983w1315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range989w1323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range995w1331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1001w1339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1007w1347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1013w1355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1019w1363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1025w1371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1031w1379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1037w1387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range875w1171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1043w1395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1049w1403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1052w1411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range850w1419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range881w1179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range887w1187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range893w1195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range899w1203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range905w1211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range911w1219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range917w1227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1720w2001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1779w2082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1785w2090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1791w2098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1797w2106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1803w2114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1809w2122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1815w2130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1821w2138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1827w2146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1833w2154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1725w2010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1839w2162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1845w2170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1851w2178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1857w2186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1863w2194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1869w2202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1875w2210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1881w2218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1887w2226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1893w2234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1731w2018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1899w2242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1902w2250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1702w2258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1705w2266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1737w2026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1743w2034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1749w2042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1755w2050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1761w2058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1767w2066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1773w2074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2571w2843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2630w2924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2636w2932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2642w2940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2648w2948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2654w2956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2660w2964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2666w2972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2672w2980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2678w2988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2684w2996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2576w2852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2690w3004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2696w3012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2702w3020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2708w3028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2714w3036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2720w3044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2726w3052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2732w3060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2738w3068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2744w3076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2582w2860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2747w3084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2549w3092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2552w3100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2554w3108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2588w2868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2594w2876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2600w2884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2606w2892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2612w2900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2618w2908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2624w2916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3417w3680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3476w3761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3482w3769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3488w3777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3494w3785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3500w3793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3506w3801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3512w3809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3518w3817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3524w3825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3530w3833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3422w3689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3536w3841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3542w3849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3548w3857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3554w3865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3560w3873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3566w3881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3572w3889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3578w3897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3584w3905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3587w3913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3428w3697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3391w3921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3394w3929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3396w3937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3398w3945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3434w3705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3440w3713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3446w3721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3452w3729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3458w3737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3464w3745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3470w3753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4258w4512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4317w4593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4323w4601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4329w4609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4335w4617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4341w4625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4347w4633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4353w4641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4359w4649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4365w4657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4371w4665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4263w4521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4377w4673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4383w4681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4389w4689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4395w4697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4401w4705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4407w4713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4413w4721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4419w4729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4422w4737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4228w4745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4269w4529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4231w4753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4233w4761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4235w4769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4237w4777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4275w4537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4281w4545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4287w4553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4293w4561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4299w4569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4305w4577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4311w4585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5094w5339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5153w5420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5159w5428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5165w5436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5171w5444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5177w5452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5183w5460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5189w5468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5195w5476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5201w5484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5207w5492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5099w5348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5213w5500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5219w5508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5225w5516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5231w5524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5237w5532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5243w5540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5249w5548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5252w5556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5060w5564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5063w5572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5105w5356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5065w5580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5067w5588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5069w5596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5071w5604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5111w5364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5117w5372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5123w5380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5129w5388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5135w5396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5141w5404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5147w5412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5925w6161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5984w6242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5990w6250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5996w6258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6002w6266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6008w6274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6014w6282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6020w6290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6026w6298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6032w6306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6038w6314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5930w6170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6044w6322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6050w6330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6056w6338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6062w6346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6068w6354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6074w6362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6077w6370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5887w6378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5890w6386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5892w6394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5936w6178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5894w6402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5896w6410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5898w6418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5900w6426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5942w6186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5948w6194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5954w6202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5960w6210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5966w6218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5972w6226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5978w6234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6751w6978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6810w7059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6816w7067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6822w7075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6828w7083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6834w7091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6840w7099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6846w7107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6852w7115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6858w7123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6864w7131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6756w6987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6870w7139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6876w7147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6882w7155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6888w7163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6894w7171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6897w7179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6709w7187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6712w7195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6714w7203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6716w7211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6762w6995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6718w7219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6720w7227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6722w7235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6724w7243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6768w7003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6774w7011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6780w7019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6786w7027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6792w7035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6798w7043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6804w7051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7715w7789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7744w7870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7747w7878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7750w7886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7753w7894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7756w7902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7759w7910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7762w7918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7765w7926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7768w7934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7771w7942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7717w7798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7774w7950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7777w7958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7780w7966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7546w7974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7549w7982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7551w7990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7553w7998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7555w8006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7557w8014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7559w8022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7720w7806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7561w8030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7563w8038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7565w8046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7567w8054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7723w7814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7726w7822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7729w7830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7732w7838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7735w7846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7738w7854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7741w7862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8525w8596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8554w8677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8557w8685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8560w8693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8563w8701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8566w8709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8569w8717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8572w8725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8575w8733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8578w8741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8581w8749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8527w8605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8584w8757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8587w8765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8360w8773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8363w8781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8365w8789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8367w8797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8369w8805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8371w8813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8373w8821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8375w8829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8530w8613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8377w8837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8379w8845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8381w8853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8383w8861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8533w8621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8536w8629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8539w8637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8542w8645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8545w8653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8548w8661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8551w8669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9330w9398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9359w9479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9362w9487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9365w9495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9368w9503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9371w9511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9374w9519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9377w9527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9380w9535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9383w9543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9386w9551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9332w9407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9389w9559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9169w9567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9172w9575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9174w9583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9176w9591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9178w9599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9180w9607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9182w9615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9184w9623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9186w9631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9335w9415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9188w9639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9190w9647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9192w9655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9194w9663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9338w9423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9341w9431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9344w9439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9347w9447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9350w9455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9353w9463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9356w9471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10130w10195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10159w10276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10162w10284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10165w10292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10168w10300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10171w10308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10174w10316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10177w10324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10180w10332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10183w10340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10186w10348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10132w10204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9973w10356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9976w10364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9978w10372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9980w10380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9982w10388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9984w10396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9986w10404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9988w10412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9990w10420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9992w10428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10135w10212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9994w10436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9996w10444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9998w10452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10000w10460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10138w10220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10141w10228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10144w10236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10147w10244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10150w10252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10153w10260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10156w10268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1055w1153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1084w1234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1087w1242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1090w1250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1093w1258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1096w1266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1099w1274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1102w1282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1105w1290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1108w1298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1111w1306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1057w1162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1114w1314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1117w1322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1120w1330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1123w1338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1126w1346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1129w1354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1132w1362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1135w1370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1138w1378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1141w1386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1060w1170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1144w1394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range854w1402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range857w1410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range859w1418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1063w1178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1066w1186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1069w1194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1072w1202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1075w1210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1078w1218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1081w1226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1905w2000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1934w2081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1937w2089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1940w2097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1943w2105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1946w2113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1949w2121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1952w2129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1955w2137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1958w2145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1961w2153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1907w2009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1964w2161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1967w2169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1970w2177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1973w2185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1976w2193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1979w2201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1982w2209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1985w2217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1988w2225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1991w2233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1910w2017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1708w2241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1711w2249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1713w2257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1715w2265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1913w2025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1916w2033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1919w2041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1922w2049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1925w2057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1928w2065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1931w2073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2750w2842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2779w2923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2782w2931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2785w2939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2788w2947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2791w2955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2794w2963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2797w2971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2800w2979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2803w2987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2806w2995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2752w2851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2809w3003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2812w3011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2815w3019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2818w3027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2821w3035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2824w3043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2827w3051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2830w3059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2833w3067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2557w3075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2755w2859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2560w3083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2562w3091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2564w3099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2566w3107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2758w2867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2761w2875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2764w2883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2767w2891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2770w2899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2773w2907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2776w2915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3590w3679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3619w3760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3622w3768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3625w3776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3628w3784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3631w3792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3634w3800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3637w3808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3640w3816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3643w3824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3646w3832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3592w3688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3649w3840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3652w3848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3655w3856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3658w3864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3661w3872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3664w3880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3667w3888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3670w3896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3401w3904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3404w3912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3595w3696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3406w3920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3408w3928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3410w3936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3412w3944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3598w3704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3601w3712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3604w3720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3607w3728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3610w3736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3613w3744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3616w3752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4425w4511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4454w4592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4457w4600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4460w4608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4463w4616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4466w4624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4469w4632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4472w4640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4475w4648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4478w4656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4481w4664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4427w4520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4484w4672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4487w4680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4490w4688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4493w4696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4496w4704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4499w4712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4502w4720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4240w4728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4243w4736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4245w4744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4430w4528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4247w4752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4249w4760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4251w4768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4253w4776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4433w4536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4436w4544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4439w4552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4442w4560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4445w4568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4448w4576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4451w4584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5255w5338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5284w5419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5287w5427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5290w5435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5293w5443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5296w5451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5299w5459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5302w5467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5305w5475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5308w5483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5311w5491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5257w5347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5314w5499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5317w5507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5320w5515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5323w5523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5326w5531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5329w5539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5074w5547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5077w5555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5079w5563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5081w5571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5260w5355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5083w5579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5085w5587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5087w5595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5089w5603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5263w5363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5266w5371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5269w5379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5272w5387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5275w5395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5278w5403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5281w5411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6080w6160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6109w6241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6112w6249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6115w6257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6118w6265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6121w6273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6124w6281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6127w6289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6130w6297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6133w6305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6136w6313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6082w6169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6139w6321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6142w6329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6145w6337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6148w6345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6151w6353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5903w6361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5906w6369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5908w6377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5910w6385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5912w6393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6085w6177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5914w6401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5916w6409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5918w6417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5920w6425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6088w6185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6091w6193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6094w6201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6097w6209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6100w6217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6103w6225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6106w6233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6900w6977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6929w7058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6932w7066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6935w7074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6938w7082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6941w7090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6944w7098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6947w7106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6950w7114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6953w7122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6956w7130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6902w6986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6959w7138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6962w7146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6965w7154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6968w7162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6727w7170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6730w7178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6732w7186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6734w7194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6736w7202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6738w7210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6905w6994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6740w7218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6742w7226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6744w7234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6746w7242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6908w7002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6911w7010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6914w7018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6917w7026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6920w7034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6923w7042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6926w7050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_indexbit412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8871w8873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8952w8954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8960w8962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8968w8970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8976w8978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8984w8986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8992w8994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9000w9002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9008w9010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9016w9018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9024w9026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8880w8882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9032w9034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9040w9042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9048w9050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9056w9058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9064w9066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9072w9074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9080w9082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9088w9090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9096w9098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9104w9106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8888w8890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9112w9114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9120w9122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9128w9130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9136w9138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8896w8898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8904w8906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8912w8914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8920w8922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8928w8930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8936w8938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8944w8946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9673w9675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9754w9756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9762w9764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9770w9772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9778w9780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9786w9788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9794w9796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9802w9804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9810w9812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9818w9820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9826w9828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9682w9684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9834w9836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9842w9844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9850w9852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9858w9860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9866w9868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9874w9876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9882w9884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9890w9892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9898w9900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9906w9908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9690w9692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9914w9916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9922w9924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9930w9932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9938w9940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9698w9700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9706w9708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9714w9716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9722w9724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9730w9732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9738w9740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9746w9748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10470w10472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10551w10553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10559w10561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10567w10569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10575w10577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10583w10585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10591w10593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10599w10601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10607w10609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10615w10617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10623w10625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10479w10481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10631w10633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10639w10641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10647w10649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10655w10657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10663w10665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10671w10673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10679w10681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10687w10689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10695w10697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10703w10705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10487w10489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10711w10713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10719w10721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10727w10729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10735w10737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10495w10497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10503w10505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10511w10513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10519w10521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10527w10529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10535w10537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10543w10545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1428w1430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1509w1511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1517w1519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1525w1527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1533w1535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1541w1543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1549w1551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1557w1559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1565w1567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1573w1575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1581w1583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1437w1439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1589w1591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1597w1599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1605w1607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1613w1615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1621w1623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1629w1631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1637w1639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1645w1647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1653w1655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1661w1663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1445w1447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1669w1671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1677w1679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1685w1687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1693w1695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1453w1455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1461w1463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1469w1471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1477w1479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1485w1487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1493w1495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1501w1503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2275w2277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2356w2358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2364w2366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2372w2374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2380w2382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2388w2390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2396w2398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2404w2406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2412w2414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2420w2422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2428w2430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2284w2286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2436w2438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2444w2446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2452w2454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2460w2462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2468w2470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2476w2478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2484w2486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2492w2494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2500w2502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2508w2510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2292w2294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2516w2518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2524w2526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2532w2534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2540w2542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2300w2302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2308w2310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2316w2318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2324w2326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2332w2334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2340w2342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2348w2350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3117w3119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3198w3200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3206w3208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3214w3216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3222w3224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3230w3232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3238w3240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3246w3248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3254w3256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3262w3264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3270w3272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3126w3128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3278w3280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3286w3288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3294w3296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3302w3304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3310w3312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3318w3320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3326w3328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3334w3336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3342w3344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3350w3352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3134w3136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3358w3360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3366w3368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3374w3376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3382w3384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3142w3144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3150w3152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3158w3160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3166w3168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3174w3176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3182w3184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3190w3192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3954w3956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4035w4037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4043w4045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4051w4053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4059w4061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4067w4069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4075w4077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4083w4085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4091w4093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4099w4101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4107w4109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3963w3965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4115w4117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4123w4125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4131w4133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4139w4141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4147w4149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4155w4157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4163w4165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4171w4173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4179w4181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4187w4189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3971w3973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4195w4197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4203w4205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4211w4213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4219w4221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3979w3981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3987w3989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3995w3997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4003w4005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4011w4013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4019w4021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4027w4029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4786w4788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4867w4869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4875w4877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4883w4885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4891w4893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4899w4901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4907w4909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4915w4917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4923w4925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4931w4933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4939w4941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4795w4797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4947w4949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4955w4957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4963w4965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4971w4973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4979w4981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4987w4989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4995w4997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5003w5005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5011w5013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5019w5021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4803w4805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5027w5029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5035w5037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5043w5045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5051w5053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4811w4813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4819w4821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4827w4829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4835w4837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4843w4845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4851w4853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4859w4861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5613w5615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5694w5696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5702w5704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5710w5712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5718w5720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5726w5728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5734w5736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5742w5744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5750w5752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5758w5760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5766w5768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5622w5624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5774w5776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5782w5784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5790w5792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5798w5800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5806w5808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5814w5816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5822w5824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5830w5832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5838w5840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5846w5848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5630w5632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5854w5856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5862w5864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5870w5872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5878w5880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5638w5640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5646w5648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5654w5656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5662w5664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5670w5672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5678w5680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5686w5688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6435w6437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6516w6518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6524w6526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6532w6534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6540w6542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6548w6550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6556w6558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6564w6566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6572w6574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6580w6582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6588w6590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6444w6446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6596w6598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6604w6606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6612w6614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6620w6622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6628w6630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6636w6638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6644w6646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6652w6654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6660w6662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6668w6670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6452w6454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6676w6678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6684w6686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6692w6694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6700w6702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6460w6462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6468w6470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6476w6478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6484w6486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6492w6494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6500w6502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6508w6510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7252w7254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7333w7335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7341w7343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7349w7351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7357w7359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7365w7367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7373w7375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7381w7383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7389w7391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7397w7399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7405w7407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7261w7263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7413w7415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7421w7423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7429w7431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7437w7439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7445w7447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7453w7455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7461w7463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7469w7471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7477w7479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7485w7487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7269w7271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7493w7495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7501w7503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7509w7511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7517w7519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7277w7279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7285w7287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7293w7295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7301w7303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7309w7311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7317w7319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7325w7327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8064w8066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8145w8147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8153w8155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8161w8163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8169w8171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8177w8179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8185w8187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8193w8195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8201w8203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8209w8211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8217w8219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8073w8075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8225w8227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8233w8235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8241w8243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8249w8251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8257w8259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8265w8267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8273w8275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8281w8283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8289w8291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8297w8299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8081w8083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8305w8307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8313w8315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8321w8323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8329w8331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8089w8091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8097w8099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8105w8107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8113w8115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8121w8123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8129w8131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8137w8139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10751w10755w10756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10794w10807w10808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10799w10812w10813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10804w10817w10818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10809w10822w10823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10814w10827w10828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10819w10832w10833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10824w10837w10838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10829w10842w10843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10834w10847w10848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10839w10852w10853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10759w10762w10763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10844w10857w10858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10849w10862w10863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10854w10867w10868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10859w10872w10873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10864w10877w10878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10869w10882w10883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10874w10887w10888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10879w10892w10893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10884w10897w10898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10889w10902w10903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10750w10767w10768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10894w10907w10908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10899w10912w10913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10904w10915w10916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10909w10918w10919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10758w10772w10773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10764w10777w10778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10769w10782w10783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10774w10787w10788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10779w10792w10793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10784w10797w10798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10789w10802w10803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range458w461w462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range463w466w467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range468w471w472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range473w476w477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range478w481w482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range483w486w487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range488w491w492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range493w496w497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range498w501w502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range503w506w507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range508w511w512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range513w516w517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range518w521w522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range523w526w527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range528w531w532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range533w536w537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range538w541w542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range543w546w547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range548w551w552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range553w556w557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range418w421w422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range558w561w562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range563w566w567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range568w571w572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range573w576w577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range423w426w427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range428w431w432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range433w436w437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range438w441w442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range443w446w447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range448w451w452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range453w456w457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7569w7785w7786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7628w7867w7868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7634w7875w7876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7640w7883w7884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7646w7891w7892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7652w7899w7900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7658w7907w7908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7664w7915w7916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7670w7923w7924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7676w7931w7932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7682w7939w7940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7574w7795w7796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7688w7947w7948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7694w7955w7956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7700w7963w7964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7706w7971w7972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7711w7979w7980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7522w7987w7988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7528w7995w7996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7530w8003w8004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7532w8011w8012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7534w8019w8020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7580w7803w7804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7536w8027w8028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7538w8035w8036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7540w8043w8044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7542w8051w8052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7586w7811w7812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7592w7819w7820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7598w7827w7828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7604w7835w7836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7610w7843w7844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7616w7851w7852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7622w7859w7860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8385w8592w8593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8444w8674w8675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8450w8682w8683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8456w8690w8691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8462w8698w8699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8468w8706w8707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8474w8714w8715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8480w8722w8723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8486w8730w8731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8492w8738w8739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8498w8746w8747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8390w8602w8603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8504w8754w8755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8510w8762w8763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8516w8770w8771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8521w8778w8779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8334w8786w8787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8340w8794w8795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8342w8802w8803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8344w8810w8811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8346w8818w8819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8348w8826w8827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8396w8610w8611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8350w8834w8835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8352w8842w8843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8354w8850w8851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8356w8858w8859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8402w8618w8619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8408w8626w8627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8414w8634w8635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8420w8642w8643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8426w8650w8651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8432w8658w8659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8438w8666w8667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9196w9394w9395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9255w9476w9477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9261w9484w9485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9267w9492w9493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9273w9500w9501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9279w9508w9509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9285w9516w9517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9291w9524w9525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9297w9532w9533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9303w9540w9541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9309w9548w9549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9201w9404w9405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9315w9556w9557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9321w9564w9565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9326w9572w9573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9141w9580w9581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9147w9588w9589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9149w9596w9597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9151w9604w9605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9153w9612w9613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9155w9620w9621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9157w9628w9629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9207w9412w9413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9159w9636w9637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9161w9644w9645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9163w9652w9653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9165w9660w9661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9213w9420w9421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9219w9428w9429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9225w9436w9437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9231w9444w9445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9237w9452w9453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9243w9460w9461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9249w9468w9469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range861w1149w1150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range920w1231w1232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range926w1239w1240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range932w1247w1248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range938w1255w1256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range944w1263w1264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range950w1271w1272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range956w1279w1280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range962w1287w1288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range968w1295w1296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range974w1303w1304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range866w1159w1160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range980w1311w1312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range986w1319w1320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range992w1327w1328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range998w1335w1336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1004w1343w1344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1010w1351w1352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1016w1359w1360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1022w1367w1368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1028w1375w1376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1034w1383w1384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range872w1167w1168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1040w1391w1392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1046w1399w1400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1051w1407w1408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range846w1415w1416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range878w1175w1176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range884w1183w1184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range890w1191w1192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range896w1199w1200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range902w1207w1208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range908w1215w1216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range914w1223w1224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1717w1996w1997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1776w2078w2079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1782w2086w2087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1788w2094w2095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1794w2102w2103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1800w2110w2111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1806w2118w2119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1812w2126w2127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1818w2134w2135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1824w2142w2143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1830w2150w2151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1722w2006w2007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1836w2158w2159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1842w2166w2167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1848w2174w2175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1854w2182w2183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1860w2190w2191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1866w2198w2199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1872w2206w2207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1878w2214w2215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1884w2222w2223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1890w2230w2231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1728w2014w2015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1896w2238w2239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1901w2246w2247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1698w2254w2255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1704w2262w2263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1734w2022w2023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1740w2030w2031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1746w2038w2039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1752w2046w2047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1758w2054w2055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1764w2062w2063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1770w2070w2071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2568w2838w2839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2627w2920w2921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2633w2928w2929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2639w2936w2937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2645w2944w2945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2651w2952w2953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2657w2960w2961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2663w2968w2969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2669w2976w2977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2675w2984w2985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2681w2992w2993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2573w2848w2849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2687w3000w3001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2693w3008w3009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2699w3016w3017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2705w3024w3025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2711w3032w3033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2717w3040w3041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2723w3048w3049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2729w3056w3057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2735w3064w3065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2741w3072w3073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2579w2856w2857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2746w3080w3081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2545w3088w3089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2551w3096w3097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2553w3104w3105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2585w2864w2865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2591w2872w2873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2597w2880w2881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2603w2888w2889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2609w2896w2897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2615w2904w2905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2621w2912w2913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3414w3675w3676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3473w3757w3758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3479w3765w3766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3485w3773w3774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3491w3781w3782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3497w3789w3790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3503w3797w3798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3509w3805w3806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3515w3813w3814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3521w3821w3822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3527w3829w3830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3419w3685w3686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3533w3837w3838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3539w3845w3846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3545w3853w3854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3551w3861w3862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3557w3869w3870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3563w3877w3878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3569w3885w3886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3575w3893w3894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3581w3901w3902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3586w3909w3910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3425w3693w3694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3387w3917w3918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3393w3925w3926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3395w3933w3934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3397w3941w3942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3431w3701w3702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3437w3709w3710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3443w3717w3718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3449w3725w3726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3455w3733w3734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3461w3741w3742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3467w3749w3750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4255w4507w4508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4314w4589w4590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4320w4597w4598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4326w4605w4606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4332w4613w4614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4338w4621w4622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4344w4629w4630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4350w4637w4638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4356w4645w4646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4362w4653w4654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4368w4661w4662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4260w4517w4518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4374w4669w4670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4380w4677w4678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4386w4685w4686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4392w4693w4694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4398w4701w4702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4404w4709w4710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4410w4717w4718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4416w4725w4726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4421w4733w4734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4224w4741w4742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4266w4525w4526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4230w4749w4750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4232w4757w4758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4234w4765w4766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4236w4773w4774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4272w4533w4534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4278w4541w4542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4284w4549w4550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4290w4557w4558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4296w4565w4566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4302w4573w4574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4308w4581w4582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5091w5334w5335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5150w5416w5417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5156w5424w5425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5162w5432w5433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5168w5440w5441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5174w5448w5449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5180w5456w5457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5186w5464w5465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5192w5472w5473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5198w5480w5481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5204w5488w5489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5096w5344w5345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5210w5496w5497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5216w5504w5505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5222w5512w5513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5228w5520w5521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5234w5528w5529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5240w5536w5537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5246w5544w5545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5251w5552w5553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5056w5560w5561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5062w5568w5569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5102w5352w5353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5064w5576w5577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5066w5584w5585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5068w5592w5593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5070w5600w5601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5108w5360w5361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5114w5368w5369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5120w5376w5377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5126w5384w5385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5132w5392w5393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5138w5400w5401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5144w5408w5409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5922w6156w6157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5981w6238w6239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5987w6246w6247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5993w6254w6255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5999w6262w6263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6005w6270w6271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6011w6278w6279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6017w6286w6287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6023w6294w6295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6029w6302w6303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6035w6310w6311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5927w6166w6167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6041w6318w6319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6047w6326w6327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6053w6334w6335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6059w6342w6343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6065w6350w6351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6071w6358w6359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6076w6366w6367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5883w6374w6375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5889w6382w6383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5891w6390w6391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5933w6174w6175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5893w6398w6399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5895w6406w6407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5897w6414w6415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5899w6422w6423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5939w6182w6183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5945w6190w6191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5951w6198w6199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5957w6206w6207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5963w6214w6215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5969w6222w6223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5975w6230w6231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6748w6973w6974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6807w7055w7056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6813w7063w7064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6819w7071w7072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6825w7079w7080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6831w7087w7088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6837w7095w7096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6843w7103w7104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6849w7111w7112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6855w7119w7120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6861w7127w7128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6753w6983w6984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6867w7135w7136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6873w7143w7144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6879w7151w7152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6885w7159w7160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6891w7167w7168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6896w7175w7176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6705w7183w7184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6711w7191w7192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6713w7199w7200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6715w7207w7208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6759w6991w6992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6717w7215w7216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6719w7223w7224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6721w7231w7232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6723w7239w7240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6765w6999w7000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6771w7007w7008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6777w7015w7016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6783w7023w7024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6789w7031w7032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6795w7039w7040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6801w7047w7048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7572w7790w7791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7631w7871w7872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7637w7879w7880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7643w7887w7888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7649w7895w7896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7655w7903w7904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7661w7911w7912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7667w7919w7920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7673w7927w7928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7679w7935w7936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7685w7943w7944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7577w7799w7800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7691w7951w7952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7697w7959w7960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7703w7967w7968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7709w7975w7976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7712w7983w7984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7526w7991w7992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7529w7999w8000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7531w8007w8008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7533w8015w8016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7535w8023w8024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7583w7807w7808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7537w8031w8032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7539w8039w8040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7541w8047w8048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7543w8055w8056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7589w7815w7816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7595w7823w7824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7601w7831w7832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7607w7839w7840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7613w7847w7848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7619w7855w7856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7625w7863w7864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8388w8597w8598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8447w8678w8679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8453w8686w8687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8459w8694w8695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8465w8702w8703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8471w8710w8711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8477w8718w8719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8483w8726w8727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8489w8734w8735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8495w8742w8743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8501w8750w8751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8393w8606w8607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8507w8758w8759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8513w8766w8767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8519w8774w8775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8522w8782w8783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8338w8790w8791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8341w8798w8799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8343w8806w8807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8345w8814w8815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8347w8822w8823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8349w8830w8831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8399w8614w8615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8351w8838w8839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8353w8846w8847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8355w8854w8855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8357w8862w8863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8405w8622w8623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8411w8630w8631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8417w8638w8639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8423w8646w8647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8429w8654w8655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8435w8662w8663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8441w8670w8671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9199w9399w9400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9258w9480w9481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9264w9488w9489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9270w9496w9497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9276w9504w9505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9282w9512w9513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9288w9520w9521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9294w9528w9529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9300w9536w9537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9306w9544w9545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9312w9552w9553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9204w9408w9409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9318w9560w9561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9324w9568w9569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9327w9576w9577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9145w9584w9585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9148w9592w9593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9150w9600w9601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9152w9608w9609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9154w9616w9617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9156w9624w9625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9158w9632w9633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9210w9416w9417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9160w9640w9641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9162w9648w9649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9164w9656w9657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9166w9664w9665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9216w9424w9425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9222w9432w9433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9228w9440w9441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9234w9448w9449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9240w9456w9457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9246w9464w9465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9252w9472w9473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range864w1154w1155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range923w1235w1236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range929w1243w1244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range935w1251w1252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range941w1259w1260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range947w1267w1268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range953w1275w1276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range959w1283w1284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range965w1291w1292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range971w1299w1300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range977w1307w1308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range869w1163w1164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range983w1315w1316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range989w1323w1324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range995w1331w1332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1001w1339w1340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1007w1347w1348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1013w1355w1356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1019w1363w1364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1025w1371w1372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1031w1379w1380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1037w1387w1388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range875w1171w1172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1043w1395w1396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1049w1403w1404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1052w1411w1412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range850w1419w1420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range881w1179w1180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range887w1187w1188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range893w1195w1196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range899w1203w1204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range905w1211w1212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range911w1219w1220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range917w1227w1228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1720w2001w2002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1779w2082w2083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1785w2090w2091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1791w2098w2099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1797w2106w2107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1803w2114w2115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1809w2122w2123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1815w2130w2131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1821w2138w2139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1827w2146w2147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1833w2154w2155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1725w2010w2011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1839w2162w2163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1845w2170w2171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1851w2178w2179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1857w2186w2187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1863w2194w2195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1869w2202w2203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1875w2210w2211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1881w2218w2219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1887w2226w2227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1893w2234w2235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1731w2018w2019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1899w2242w2243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1902w2250w2251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1702w2258w2259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1705w2266w2267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1737w2026w2027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1743w2034w2035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1749w2042w2043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1755w2050w2051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1761w2058w2059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1767w2066w2067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1773w2074w2075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2571w2843w2844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2630w2924w2925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2636w2932w2933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2642w2940w2941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2648w2948w2949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2654w2956w2957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2660w2964w2965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2666w2972w2973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2672w2980w2981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2678w2988w2989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2684w2996w2997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2576w2852w2853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2690w3004w3005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2696w3012w3013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2702w3020w3021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2708w3028w3029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2714w3036w3037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2720w3044w3045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2726w3052w3053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2732w3060w3061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2738w3068w3069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2744w3076w3077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2582w2860w2861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2747w3084w3085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2549w3092w3093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2552w3100w3101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2554w3108w3109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2588w2868w2869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2594w2876w2877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2600w2884w2885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2606w2892w2893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2612w2900w2901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2618w2908w2909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2624w2916w2917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3417w3680w3681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3476w3761w3762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3482w3769w3770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3488w3777w3778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3494w3785w3786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3500w3793w3794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3506w3801w3802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3512w3809w3810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3518w3817w3818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3524w3825w3826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3530w3833w3834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3422w3689w3690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3536w3841w3842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3542w3849w3850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3548w3857w3858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3554w3865w3866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3560w3873w3874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3566w3881w3882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3572w3889w3890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3578w3897w3898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3584w3905w3906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3587w3913w3914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3428w3697w3698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3391w3921w3922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3394w3929w3930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3396w3937w3938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3398w3945w3946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3434w3705w3706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3440w3713w3714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3446w3721w3722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3452w3729w3730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3458w3737w3738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3464w3745w3746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3470w3753w3754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4258w4512w4513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4317w4593w4594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4323w4601w4602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4329w4609w4610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4335w4617w4618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4341w4625w4626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4347w4633w4634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4353w4641w4642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4359w4649w4650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4365w4657w4658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4371w4665w4666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4263w4521w4522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4377w4673w4674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4383w4681w4682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4389w4689w4690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4395w4697w4698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4401w4705w4706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4407w4713w4714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4413w4721w4722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4419w4729w4730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4422w4737w4738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4228w4745w4746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4269w4529w4530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4231w4753w4754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4233w4761w4762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4235w4769w4770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4237w4777w4778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4275w4537w4538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4281w4545w4546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4287w4553w4554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4293w4561w4562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4299w4569w4570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4305w4577w4578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4311w4585w4586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5094w5339w5340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5153w5420w5421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5159w5428w5429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5165w5436w5437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5171w5444w5445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5177w5452w5453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5183w5460w5461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5189w5468w5469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5195w5476w5477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5201w5484w5485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5207w5492w5493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5099w5348w5349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5213w5500w5501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5219w5508w5509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5225w5516w5517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5231w5524w5525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5237w5532w5533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5243w5540w5541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5249w5548w5549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5252w5556w5557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5060w5564w5565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5063w5572w5573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5105w5356w5357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5065w5580w5581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5067w5588w5589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5069w5596w5597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5071w5604w5605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5111w5364w5365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5117w5372w5373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5123w5380w5381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5129w5388w5389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5135w5396w5397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5141w5404w5405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5147w5412w5413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5925w6161w6162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5984w6242w6243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5990w6250w6251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5996w6258w6259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6002w6266w6267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6008w6274w6275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6014w6282w6283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6020w6290w6291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6026w6298w6299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6032w6306w6307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6038w6314w6315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5930w6170w6171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6044w6322w6323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6050w6330w6331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6056w6338w6339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6062w6346w6347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6068w6354w6355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6074w6362w6363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6077w6370w6371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5887w6378w6379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5890w6386w6387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5892w6394w6395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5936w6178w6179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5894w6402w6403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5896w6410w6411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5898w6418w6419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5900w6426w6427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5942w6186w6187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5948w6194w6195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5954w6202w6203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5960w6210w6211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5966w6218w6219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5972w6226w6227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5978w6234w6235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6751w6978w6979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6810w7059w7060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6816w7067w7068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6822w7075w7076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6828w7083w7084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6834w7091w7092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6840w7099w7100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6846w7107w7108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6852w7115w7116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6858w7123w7124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6864w7131w7132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6756w6987w6988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6870w7139w7140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6876w7147w7148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6882w7155w7156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6888w7163w7164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6894w7171w7172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6897w7179w7180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6709w7187w7188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6712w7195w7196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6714w7203w7204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6716w7211w7212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6762w6995w6996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6718w7219w7220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6720w7227w7228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6722w7235w7236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6724w7243w7244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6768w7003w7004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6774w7011w7012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6780w7019w7020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6786w7027w7028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6792w7035w7036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6798w7043w7044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6804w7051w7052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8871w8873w8874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8952w8954w8955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8960w8962w8963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8968w8970w8971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8976w8978w8979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8984w8986w8987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8992w8994w8995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9000w9002w9003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9008w9010w9011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9016w9018w9019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9024w9026w9027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8880w8882w8883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9032w9034w9035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9040w9042w9043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9048w9050w9051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9056w9058w9059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9064w9066w9067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9072w9074w9075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9080w9082w9083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9088w9090w9091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9096w9098w9099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9104w9106w9107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8888w8890w8891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9112w9114w9115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9120w9122w9123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9128w9130w9131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9136w9138w9139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8896w8898w8899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8904w8906w8907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8912w8914w8915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8920w8922w8923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8928w8930w8931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8936w8938w8939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8944w8946w8947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9673w9675w9676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9754w9756w9757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9762w9764w9765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9770w9772w9773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9778w9780w9781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9786w9788w9789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9794w9796w9797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9802w9804w9805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9810w9812w9813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9818w9820w9821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9826w9828w9829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9682w9684w9685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9834w9836w9837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9842w9844w9845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9850w9852w9853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9858w9860w9861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9866w9868w9869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9874w9876w9877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9882w9884w9885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9890w9892w9893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9898w9900w9901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9906w9908w9909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9690w9692w9693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9914w9916w9917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9922w9924w9925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9930w9932w9933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9938w9940w9941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9698w9700w9701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9706w9708w9709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9714w9716w9717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9722w9724w9725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9730w9732w9733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9738w9740w9741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9746w9748w9749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10470w10472w10473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10551w10553w10554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10559w10561w10562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10567w10569w10570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10575w10577w10578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10583w10585w10586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10591w10593w10594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10599w10601w10602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10607w10609w10610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10615w10617w10618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10623w10625w10626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10479w10481w10482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10631w10633w10634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10639w10641w10642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10647w10649w10650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10655w10657w10658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10663w10665w10666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10671w10673w10674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10679w10681w10682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10687w10689w10690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10695w10697w10698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10703w10705w10706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10487w10489w10490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10711w10713w10714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10719w10721w10722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10727w10729w10730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10735w10737w10738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10495w10497w10498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10503w10505w10506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10511w10513w10514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10519w10521w10522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10527w10529w10530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10535w10537w10538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10543w10545w10546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1428w1430w1431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1509w1511w1512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1517w1519w1520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1525w1527w1528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1533w1535w1536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1541w1543w1544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1549w1551w1552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1557w1559w1560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1565w1567w1568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1573w1575w1576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1581w1583w1584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1437w1439w1440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1589w1591w1592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1597w1599w1600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1605w1607w1608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1613w1615w1616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1621w1623w1624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1629w1631w1632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1637w1639w1640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1645w1647w1648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1653w1655w1656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1661w1663w1664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1445w1447w1448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1669w1671w1672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1677w1679w1680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1685w1687w1688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1693w1695w1696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1453w1455w1456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1461w1463w1464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1469w1471w1472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1477w1479w1480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1485w1487w1488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1493w1495w1496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1501w1503w1504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2275w2277w2278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2356w2358w2359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2364w2366w2367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2372w2374w2375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2380w2382w2383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2388w2390w2391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2396w2398w2399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2404w2406w2407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2412w2414w2415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2420w2422w2423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2428w2430w2431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2284w2286w2287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2436w2438w2439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2444w2446w2447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2452w2454w2455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2460w2462w2463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2468w2470w2471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2476w2478w2479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2484w2486w2487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2492w2494w2495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2500w2502w2503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2508w2510w2511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2292w2294w2295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2516w2518w2519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2524w2526w2527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2532w2534w2535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2540w2542w2543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2300w2302w2303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2308w2310w2311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2316w2318w2319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2324w2326w2327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2332w2334w2335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2340w2342w2343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2348w2350w2351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3117w3119w3120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3198w3200w3201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3206w3208w3209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3214w3216w3217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3222w3224w3225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3230w3232w3233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3238w3240w3241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3246w3248w3249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3254w3256w3257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3262w3264w3265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3270w3272w3273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3126w3128w3129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3278w3280w3281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3286w3288w3289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3294w3296w3297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3302w3304w3305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3310w3312w3313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3318w3320w3321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3326w3328w3329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3334w3336w3337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3342w3344w3345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3350w3352w3353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3134w3136w3137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3358w3360w3361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3366w3368w3369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3374w3376w3377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3382w3384w3385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3142w3144w3145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3150w3152w3153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3158w3160w3161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3166w3168w3169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3174w3176w3177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3182w3184w3185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3190w3192w3193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3954w3956w3957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4035w4037w4038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4043w4045w4046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4051w4053w4054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4059w4061w4062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4067w4069w4070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4075w4077w4078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4083w4085w4086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4091w4093w4094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4099w4101w4102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4107w4109w4110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3963w3965w3966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4115w4117w4118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4123w4125w4126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4131w4133w4134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4139w4141w4142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4147w4149w4150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4155w4157w4158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4163w4165w4166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4171w4173w4174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4179w4181w4182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4187w4189w4190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3971w3973w3974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4195w4197w4198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4203w4205w4206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4211w4213w4214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4219w4221w4222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3979w3981w3982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3987w3989w3990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3995w3997w3998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4003w4005w4006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4011w4013w4014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4019w4021w4022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4027w4029w4030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4786w4788w4789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4867w4869w4870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4875w4877w4878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4883w4885w4886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4891w4893w4894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4899w4901w4902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4907w4909w4910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4915w4917w4918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4923w4925w4926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4931w4933w4934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4939w4941w4942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4795w4797w4798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4947w4949w4950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4955w4957w4958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4963w4965w4966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4971w4973w4974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4979w4981w4982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4987w4989w4990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4995w4997w4998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5003w5005w5006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5011w5013w5014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5019w5021w5022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4803w4805w4806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5027w5029w5030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5035w5037w5038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5043w5045w5046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5051w5053w5054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4811w4813w4814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4819w4821w4822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4827w4829w4830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4835w4837w4838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4843w4845w4846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4851w4853w4854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4859w4861w4862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5613w5615w5616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5694w5696w5697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5702w5704w5705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5710w5712w5713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5718w5720w5721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5726w5728w5729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5734w5736w5737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5742w5744w5745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5750w5752w5753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5758w5760w5761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5766w5768w5769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5622w5624w5625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5774w5776w5777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5782w5784w5785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5790w5792w5793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5798w5800w5801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5806w5808w5809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5814w5816w5817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5822w5824w5825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5830w5832w5833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5838w5840w5841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5846w5848w5849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5630w5632w5633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5854w5856w5857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5862w5864w5865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5870w5872w5873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5878w5880w5881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5638w5640w5641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5646w5648w5649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5654w5656w5657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5662w5664w5665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5670w5672w5673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5678w5680w5681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5686w5688w5689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6435w6437w6438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6516w6518w6519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6524w6526w6527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6532w6534w6535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6540w6542w6543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6548w6550w6551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6556w6558w6559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6564w6566w6567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6572w6574w6575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6580w6582w6583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6588w6590w6591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6444w6446w6447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6596w6598w6599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6604w6606w6607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6612w6614w6615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6620w6622w6623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6628w6630w6631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6636w6638w6639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6644w6646w6647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6652w6654w6655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6660w6662w6663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6668w6670w6671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6452w6454w6455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6676w6678w6679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6684w6686w6687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6692w6694w6695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6700w6702w6703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6460w6462w6463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6468w6470w6471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6476w6478w6479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6484w6486w6487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6492w6494w6495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6500w6502w6503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6508w6510w6511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7252w7254w7255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7333w7335w7336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7341w7343w7344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7349w7351w7352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7357w7359w7360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7365w7367w7368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7373w7375w7376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7381w7383w7384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7389w7391w7392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7397w7399w7400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7405w7407w7408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7261w7263w7264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7413w7415w7416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7421w7423w7424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7429w7431w7432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7437w7439w7440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7445w7447w7448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7453w7455w7456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7461w7463w7464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7469w7471w7472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7477w7479w7480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7485w7487w7488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7269w7271w7272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7493w7495w7496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7501w7503w7504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7509w7511w7512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7517w7519w7520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7277w7279w7280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7285w7287w7288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7293w7295w7296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7301w7303w7304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7309w7311w7312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7317w7319w7320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7325w7327w7328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8064w8066w8067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8145w8147w8148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8153w8155w8156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8161w8163w8164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8169w8171w8172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8177w8179w8180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8185w8187w8188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8193w8195w8196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8201w8203w8204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8209w8211w8212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8217w8219w8220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8073w8075w8076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8225w8227w8228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8233w8235w8236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8241w8243w8244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8249w8251w8252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8257w8259w8260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8265w8267w8268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8273w8275w8276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8281w8283w8284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8289w8291w8292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8297w8299w8300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8081w8083w8084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8305w8307w8308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8313w8315w8316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8321w8323w8324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8329w8331w8332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8089w8091w8092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8097w8099w8100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8105w8107w8108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8113w8115w8116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8121w8123w8124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8129w8131w8132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8137w8139w8140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_estimate_w10920w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7782w8059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7865w8142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7873w8150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7881w8158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7889w8166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7897w8174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7905w8182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7913w8190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7921w8198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7929w8206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7937w8214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7793w8070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7945w8222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7953w8230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7961w8238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7969w8246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7977w8254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7985w8262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7993w8270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8001w8278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8009w8286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8017w8294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7801w8078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8025w8302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8033w8310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8041w8318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8049w8326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7809w8086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7817w8094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7825w8102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7833w8110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7841w8118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7849w8126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7857w8134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8589w8866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8672w8949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8680w8957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8688w8965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8696w8973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8704w8981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8712w8989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8720w8997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8728w9005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8736w9013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8744w9021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8600w8877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8752w9029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8760w9037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8768w9045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8776w9053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8784w9061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8792w9069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8800w9077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8808w9085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8816w9093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8824w9101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8608w8885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8832w9109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8840w9117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8848w9125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8856w9133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8616w8893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8624w8901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8632w8909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8640w8917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8648w8925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8656w8933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8664w8941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9391w9668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9474w9751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9482w9759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9490w9767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9498w9775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9506w9783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9514w9791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9522w9799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9530w9807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9538w9815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9546w9823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9402w9679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9554w9831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9562w9839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9570w9847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9578w9855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9586w9863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9594w9871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9602w9879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9610w9887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9618w9895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9626w9903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9410w9687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9634w9911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9642w9919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9650w9927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9658w9935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9418w9695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9426w9703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9434w9711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9442w9719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9450w9727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9458w9735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9466w9743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10188w10465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10271w10548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10279w10556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10287w10564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10295w10572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10303w10580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10311w10588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10319w10596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10327w10604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10335w10612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10343w10620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10199w10476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10351w10628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10359w10636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10367w10644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10375w10652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10383w10660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10391w10668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10399w10676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10407w10684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10415w10692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10423w10700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10207w10484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10431w10708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10439w10716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10447w10724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10455w10732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10215w10492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10223w10500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10231w10508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10239w10516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10247w10524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10255w10532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10263w10540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1146w1423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1229w1506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1237w1514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1245w1522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1253w1530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1261w1538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1269w1546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1277w1554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1285w1562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1293w1570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1301w1578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1157w1434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1309w1586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1317w1594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1325w1602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1333w1610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1341w1618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1349w1626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1357w1634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1365w1642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1373w1650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1381w1658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1165w1442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1389w1666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1397w1674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1405w1682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1413w1690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1173w1450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1181w1458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1189w1466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1197w1474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1205w1482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1213w1490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1221w1498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1993w2270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2076w2353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2084w2361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2092w2369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2100w2377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2108w2385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2116w2393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2124w2401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2132w2409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2140w2417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2148w2425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2004w2281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2156w2433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2164w2441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2172w2449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2180w2457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2188w2465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2196w2473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2204w2481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2212w2489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2220w2497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2228w2505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2012w2289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2236w2513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2244w2521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2252w2529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2260w2537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2020w2297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2028w2305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2036w2313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2044w2321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2052w2329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2060w2337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2068w2345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2835w3112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2918w3195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2926w3203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2934w3211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2942w3219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2950w3227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2958w3235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2966w3243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2974w3251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2982w3259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2990w3267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2846w3123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2998w3275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3006w3283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3014w3291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3022w3299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3030w3307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3038w3315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3046w3323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3054w3331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3062w3339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3070w3347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2854w3131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3078w3355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3086w3363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3094w3371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3102w3379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2862w3139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2870w3147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2878w3155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2886w3163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2894w3171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2902w3179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2910w3187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3672w3949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3755w4032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3763w4040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3771w4048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3779w4056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3787w4064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3795w4072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3803w4080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3811w4088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3819w4096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3827w4104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3683w3960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3835w4112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3843w4120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3851w4128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3859w4136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3867w4144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3875w4152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3883w4160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3891w4168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3899w4176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3907w4184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3691w3968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3915w4192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3923w4200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3931w4208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3939w4216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3699w3976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3707w3984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3715w3992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3723w4000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3731w4008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3739w4016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3747w4024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4504w4781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4587w4864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4595w4872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4603w4880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4611w4888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4619w4896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4627w4904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4635w4912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4643w4920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4651w4928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4659w4936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4515w4792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4667w4944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4675w4952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4683w4960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4691w4968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4699w4976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4707w4984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4715w4992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4723w5000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4731w5008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4739w5016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4523w4800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4747w5024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4755w5032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4763w5040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4771w5048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4531w4808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4539w4816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4547w4824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4555w4832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4563w4840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4571w4848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4579w4856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5331w5608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5414w5691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5422w5699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5430w5707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5438w5715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5446w5723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5454w5731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5462w5739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5470w5747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5478w5755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5486w5763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5342w5619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5494w5771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5502w5779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5510w5787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5518w5795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5526w5803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5534w5811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5542w5819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5550w5827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5558w5835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5566w5843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5350w5627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5574w5851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5582w5859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5590w5867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5598w5875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5358w5635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5366w5643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5374w5651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5382w5659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5390w5667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5398w5675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5406w5683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6153w6430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6236w6513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6244w6521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6252w6529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6260w6537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6268w6545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6276w6553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6284w6561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6292w6569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6300w6577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6308w6585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6164w6441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6316w6593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6324w6601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6332w6609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6340w6617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6348w6625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6356w6633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6364w6641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6372w6649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6380w6657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6388w6665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6172w6449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6396w6673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6404w6681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6412w6689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6420w6697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6180w6457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6188w6465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6196w6473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6204w6481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6212w6489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6220w6497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6228w6505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6970w7247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7053w7330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7061w7338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7069w7346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7077w7354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7085w7362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7093w7370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7101w7378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7109w7386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7117w7394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7125w7402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6981w7258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7133w7410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7141w7418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7149w7426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7157w7434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7165w7442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7173w7450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7181w7458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7189w7466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7197w7474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7205w7482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6989w7266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7213w7490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7221w7498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7229w7506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7237w7514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6997w7274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7005w7282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7013w7290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7021w7298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7029w7306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7037w7314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7045w7322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7788w8062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7869w8144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7877w8152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7885w8160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7893w8168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7901w8176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7909w8184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7917w8192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7925w8200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7933w8208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7941w8216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7797w8072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7949w8224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7957w8232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7965w8240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7973w8248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7981w8256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7989w8264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7997w8272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8005w8280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8013w8288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8021w8296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7805w8080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8029w8304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8037w8312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8045w8320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8053w8328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7813w8088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7821w8096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7829w8104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7837w8112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7845w8120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7853w8128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7861w8136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8595w8869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8676w8951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8684w8959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8692w8967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8700w8975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8708w8983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8716w8991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8724w8999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8732w9007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8740w9015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8748w9023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8604w8879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8756w9031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8764w9039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8772w9047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8780w9055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8788w9063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8796w9071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8804w9079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8812w9087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8820w9095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8828w9103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8612w8887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8836w9111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8844w9119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8852w9127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8860w9135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8620w8895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8628w8903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8636w8911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8644w8919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8652w8927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8660w8935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8668w8943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9397w9671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9478w9753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9486w9761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9494w9769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9502w9777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9510w9785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9518w9793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9526w9801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9534w9809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9542w9817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9550w9825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9406w9681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9558w9833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9566w9841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9574w9849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9582w9857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9590w9865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9598w9873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9606w9881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9614w9889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9622w9897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9630w9905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9414w9689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9638w9913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9646w9921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9654w9929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9662w9937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9422w9697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9430w9705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9438w9713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9446w9721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9454w9729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9462w9737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9470w9745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10194w10468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10275w10550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10283w10558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10291w10566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10299w10574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10307w10582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10315w10590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10323w10598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10331w10606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10339w10614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10347w10622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10203w10478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10355w10630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10363w10638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10371w10646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10379w10654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10387w10662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10395w10670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10403w10678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10411w10686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10419w10694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10427w10702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10211w10486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10435w10710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10443w10718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10451w10726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10459w10734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10219w10494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10227w10502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10235w10510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10243w10518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10251w10526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10259w10534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10267w10542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1152w1426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1233w1508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1241w1516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1249w1524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1257w1532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1265w1540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1273w1548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1281w1556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1289w1564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1297w1572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1305w1580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1161w1436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1313w1588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1321w1596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1329w1604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1337w1612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1345w1620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1353w1628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1361w1636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1369w1644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1377w1652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1385w1660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1169w1444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1393w1668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1401w1676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1409w1684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1417w1692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1177w1452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1185w1460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1193w1468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1201w1476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1209w1484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1217w1492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1225w1500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1999w2273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2080w2355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2088w2363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2096w2371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2104w2379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2112w2387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2120w2395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2128w2403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2136w2411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2144w2419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2152w2427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2008w2283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2160w2435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2168w2443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2176w2451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2184w2459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2192w2467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2200w2475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2208w2483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2216w2491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2224w2499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2232w2507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2016w2291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2240w2515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2248w2523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2256w2531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2264w2539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2024w2299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2032w2307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2040w2315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2048w2323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2056w2331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2064w2339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2072w2347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2841w3115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2922w3197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2930w3205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2938w3213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2946w3221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2954w3229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2962w3237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2970w3245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2978w3253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2986w3261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2994w3269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2850w3125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3002w3277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3010w3285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3018w3293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3026w3301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3034w3309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3042w3317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3050w3325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3058w3333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3066w3341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3074w3349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2858w3133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3082w3357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3090w3365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3098w3373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3106w3381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2866w3141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2874w3149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2882w3157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2890w3165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2898w3173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2906w3181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2914w3189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3678w3952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3759w4034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3767w4042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3775w4050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3783w4058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3791w4066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3799w4074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3807w4082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3815w4090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3823w4098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3831w4106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3687w3962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3839w4114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3847w4122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3855w4130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3863w4138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3871w4146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3879w4154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3887w4162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3895w4170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3903w4178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3911w4186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3695w3970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3919w4194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3927w4202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3935w4210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3943w4218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3703w3978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3711w3986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3719w3994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3727w4002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3735w4010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3743w4018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3751w4026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4510w4784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4591w4866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4599w4874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4607w4882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4615w4890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4623w4898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4631w4906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4639w4914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4647w4922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4655w4930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4663w4938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4519w4794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4671w4946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4679w4954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4687w4962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4695w4970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4703w4978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4711w4986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4719w4994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4727w5002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4735w5010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4743w5018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4527w4802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4751w5026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4759w5034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4767w5042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4775w5050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4535w4810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4543w4818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4551w4826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4559w4834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4567w4842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4575w4850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4583w4858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5337w5611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5418w5693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5426w5701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5434w5709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5442w5717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5450w5725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5458w5733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5466w5741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5474w5749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5482w5757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5490w5765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5346w5621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5498w5773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5506w5781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5514w5789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5522w5797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5530w5805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5538w5813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5546w5821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5554w5829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5562w5837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5570w5845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5354w5629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5578w5853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5586w5861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5594w5869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5602w5877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5362w5637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5370w5645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5378w5653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5386w5661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5394w5669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5402w5677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5410w5685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6159w6433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6240w6515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6248w6523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6256w6531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6264w6539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6272w6547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6280w6555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6288w6563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6296w6571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6304w6579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6312w6587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6168w6443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6320w6595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6328w6603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6336w6611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6344w6619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6352w6627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6360w6635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6368w6643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6376w6651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6384w6659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6392w6667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6176w6451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6400w6675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6408w6683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6416w6691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6424w6699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6184w6459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6192w6467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6200w6475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6208w6483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6216w6491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6224w6499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6232w6507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6976w7250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7057w7332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7065w7340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7073w7348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7081w7356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7089w7364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7097w7372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7105w7380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7113w7388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7121w7396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7129w7404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6985w7260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7137w7412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7145w7420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7153w7428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7161w7436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7169w7444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7177w7452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7185w7460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7193w7468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7201w7476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7209w7484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6993w7268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7217w7492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7225w7500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7233w7508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7241w7516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7001w7276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7009w7284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7017w7292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7025w7300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7033w7308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7041w7316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7049w7324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  atannode_0_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_1_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  delay_input_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  delay_pipe_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  estimate_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  indexpointnum_w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  multiplier_input_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  multipliernode_w :	STD_LOGIC_VECTOR (67 DOWNTO 0);
	 SIGNAL  post_estimate_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  pre_estimate_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  radians_load_node_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  startindex_w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  x_pipenode_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_pipenode_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_pipenode_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_pipenode_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_pipenode_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_pipenode_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_pipenode_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_pipenode_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_pipenode_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_pipenode_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_pipenode_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_pipenode_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_start_node_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_1_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range5003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range5011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range5019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range5027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range5035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range5043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range5051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range8001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range8009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range8017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range8025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range8033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range8041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range8049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range1004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range1010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range1016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range1022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range1028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range1034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range1040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range1046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range1051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range8005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range8013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range8021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range8029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range8037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range8045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range8053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range1001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range1007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range1013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range1019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range1025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range1031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range1037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range1043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range1049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range1052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  mysincos_altfp_sincos_cordic_atan_08b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  mysincos_altfp_sincos_cordic_atan_h9b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  mysincos_altfp_sincos_cordic_atan_i9b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  mysincos_altfp_sincos_cordic_atan_j9b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  mysincos_altfp_sincos_cordic_atan_k9b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  mysincos_altfp_sincos_cordic_atan_18b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  mysincos_altfp_sincos_cordic_atan_28b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  mysincos_altfp_sincos_cordic_atan_38b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  mysincos_altfp_sincos_cordic_atan_48b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  mysincos_altfp_sincos_cordic_atan_58b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  mysincos_altfp_sincos_cordic_atan_68b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  mysincos_altfp_sincos_cordic_atan_78b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  mysincos_altfp_sincos_cordic_atan_88b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  mysincos_altfp_sincos_cordic_atan_98b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  mysincos_altfp_sincos_cordic_start_339
	 PORT
	 ( 
		index	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		value	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_mult
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTHA	:	NATURAL;
		LPM_WIDTHB	:	NATURAL;
		LPM_WIDTHP	:	NATURAL;
		LPM_WIDTHS	:	NATURAL := 1;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_mult"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTHA-1 DOWNTO 0);
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTHB-1 DOWNTO 0);
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHP-1 DOWNTO 0);
		sum	:	IN STD_LOGIC_VECTOR(LPM_WIDTHS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	loop30 : FOR i IN 0 TO 3 GENERATE 
		wire_ccc_cordic_m_w_lg_indexpointnum_w409w(i) <= indexpointnum_w(i) AND indexbit;
	END GENERATE loop30;
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10751w10755w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10751w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10794w10807w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10794w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10794w10796w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10794w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10799w10812w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10799w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10799w10801w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10799w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10804w10817w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10804w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10804w10806w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10804w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10809w10822w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10809w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10809w10811w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10809w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10814w10827w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10814w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10814w10816w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10814w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10819w10832w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10819w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10819w10821w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10819w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10824w10837w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10824w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10824w10826w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10824w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10829w10842w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10829w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10829w10831w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10829w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10834w10847w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10834w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10834w10836w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10834w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10839w10852w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10839w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10839w10841w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10839w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10759w10762w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10759w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10844w10857w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10844w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10844w10846w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10844w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10849w10862w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10849w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10849w10851w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10849w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10854w10867w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10854w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10854w10856w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10854w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10859w10872w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10859w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10859w10861w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10859w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10864w10877w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10864w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10864w10866w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10864w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10869w10882w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10869w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10869w10871w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10869w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10874w10887w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10874w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10874w10876w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10874w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10879w10892w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10879w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10879w10881w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10879w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10884w10897w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10884w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10884w10886w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10884w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10889w10902w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10889w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10889w10891w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10889w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10750w10767w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10750w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10750w10753w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10750w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10894w10907w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10894w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10894w10896w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10894w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10899w10912w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10899w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10899w10901w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10899w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10904w10915w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10904w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10904w10906w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10904w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10909w10918w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10909w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10909w10911w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10909w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10758w10772w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10758w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10758w10761w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10758w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10764w10777w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10764w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10764w10766w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10764w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10769w10782w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10769w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10769w10771w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10769w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10774w10787w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10774w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10774w10776w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10774w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10779w10792w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10779w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10779w10781w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10779w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10784w10797w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10784w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10784w10786w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10784w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10789w10802w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10789w(0) AND wire_indexbitff_w_lg_w_q_range10749w10754w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10789w10791w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10789w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range410w413w(0) <= wire_ccc_cordic_m_w_radians_range410w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range410w420w(0) <= wire_ccc_cordic_m_w_radians_range410w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range458w461w(0) <= wire_ccc_cordic_m_w_radians_range458w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range458w470w(0) <= wire_ccc_cordic_m_w_radians_range458w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range463w466w(0) <= wire_ccc_cordic_m_w_radians_range463w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range463w475w(0) <= wire_ccc_cordic_m_w_radians_range463w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range468w471w(0) <= wire_ccc_cordic_m_w_radians_range468w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range468w480w(0) <= wire_ccc_cordic_m_w_radians_range468w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range473w476w(0) <= wire_ccc_cordic_m_w_radians_range473w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range473w485w(0) <= wire_ccc_cordic_m_w_radians_range473w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range478w481w(0) <= wire_ccc_cordic_m_w_radians_range478w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range478w490w(0) <= wire_ccc_cordic_m_w_radians_range478w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range483w486w(0) <= wire_ccc_cordic_m_w_radians_range483w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range483w495w(0) <= wire_ccc_cordic_m_w_radians_range483w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range488w491w(0) <= wire_ccc_cordic_m_w_radians_range488w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range488w500w(0) <= wire_ccc_cordic_m_w_radians_range488w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range493w496w(0) <= wire_ccc_cordic_m_w_radians_range493w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range493w505w(0) <= wire_ccc_cordic_m_w_radians_range493w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range498w501w(0) <= wire_ccc_cordic_m_w_radians_range498w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range498w510w(0) <= wire_ccc_cordic_m_w_radians_range498w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range503w506w(0) <= wire_ccc_cordic_m_w_radians_range503w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range503w515w(0) <= wire_ccc_cordic_m_w_radians_range503w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range415w417w(0) <= wire_ccc_cordic_m_w_radians_range415w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range415w425w(0) <= wire_ccc_cordic_m_w_radians_range415w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range508w511w(0) <= wire_ccc_cordic_m_w_radians_range508w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range508w520w(0) <= wire_ccc_cordic_m_w_radians_range508w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range513w516w(0) <= wire_ccc_cordic_m_w_radians_range513w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range513w525w(0) <= wire_ccc_cordic_m_w_radians_range513w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range518w521w(0) <= wire_ccc_cordic_m_w_radians_range518w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range518w530w(0) <= wire_ccc_cordic_m_w_radians_range518w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range523w526w(0) <= wire_ccc_cordic_m_w_radians_range523w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range523w535w(0) <= wire_ccc_cordic_m_w_radians_range523w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range528w531w(0) <= wire_ccc_cordic_m_w_radians_range528w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range528w540w(0) <= wire_ccc_cordic_m_w_radians_range528w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range533w536w(0) <= wire_ccc_cordic_m_w_radians_range533w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range533w545w(0) <= wire_ccc_cordic_m_w_radians_range533w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range538w541w(0) <= wire_ccc_cordic_m_w_radians_range538w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range538w550w(0) <= wire_ccc_cordic_m_w_radians_range538w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range543w546w(0) <= wire_ccc_cordic_m_w_radians_range543w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range543w555w(0) <= wire_ccc_cordic_m_w_radians_range543w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range548w551w(0) <= wire_ccc_cordic_m_w_radians_range548w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range548w560w(0) <= wire_ccc_cordic_m_w_radians_range548w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range553w556w(0) <= wire_ccc_cordic_m_w_radians_range553w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range553w565w(0) <= wire_ccc_cordic_m_w_radians_range553w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range418w421w(0) <= wire_ccc_cordic_m_w_radians_range418w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range418w430w(0) <= wire_ccc_cordic_m_w_radians_range418w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range558w561w(0) <= wire_ccc_cordic_m_w_radians_range558w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range558w570w(0) <= wire_ccc_cordic_m_w_radians_range558w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range563w566w(0) <= wire_ccc_cordic_m_w_radians_range563w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range563w575w(0) <= wire_ccc_cordic_m_w_radians_range563w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range568w571w(0) <= wire_ccc_cordic_m_w_radians_range568w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range573w576w(0) <= wire_ccc_cordic_m_w_radians_range573w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range423w426w(0) <= wire_ccc_cordic_m_w_radians_range423w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range423w435w(0) <= wire_ccc_cordic_m_w_radians_range423w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range428w431w(0) <= wire_ccc_cordic_m_w_radians_range428w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range428w440w(0) <= wire_ccc_cordic_m_w_radians_range428w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range433w436w(0) <= wire_ccc_cordic_m_w_radians_range433w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range433w445w(0) <= wire_ccc_cordic_m_w_radians_range433w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range438w441w(0) <= wire_ccc_cordic_m_w_radians_range438w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range438w450w(0) <= wire_ccc_cordic_m_w_radians_range438w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range443w446w(0) <= wire_ccc_cordic_m_w_radians_range443w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range443w455w(0) <= wire_ccc_cordic_m_w_radians_range443w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range448w451w(0) <= wire_ccc_cordic_m_w_radians_range448w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range448w460w(0) <= wire_ccc_cordic_m_w_radians_range448w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range453w456w(0) <= wire_ccc_cordic_m_w_radians_range453w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range453w465w(0) <= wire_ccc_cordic_m_w_radians_range453w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7569w7785w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7569w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7628w7867w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7628w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7634w7875w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7634w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7640w7883w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7640w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7646w7891w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7646w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7652w7899w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7652w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7658w7907w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7658w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7664w7915w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7664w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7670w7923w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7670w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7676w7931w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7676w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7682w7939w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7682w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7574w7795w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7574w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7688w7947w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7688w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7694w7955w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7694w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7700w7963w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7700w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7706w7971w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7706w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7711w7979w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7711w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7522w7987w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7522w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7528w7995w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7528w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7530w8003w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7530w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7532w8011w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7532w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7534w8019w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7534w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7580w7803w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7580w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7536w8027w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7536w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7538w8035w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7538w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7540w8043w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7540w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7542w8051w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7542w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7586w7811w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7586w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7592w7819w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7592w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7598w7827w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7598w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7604w7835w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7604w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7610w7843w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7610w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7616w7851w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7616w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7622w7859w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7622w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8385w8592w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8385w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8444w8674w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8444w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8450w8682w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8450w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8456w8690w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8456w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8462w8698w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8462w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8468w8706w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8468w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8474w8714w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8474w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8480w8722w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8480w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8486w8730w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8486w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8492w8738w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8492w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8498w8746w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8498w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8390w8602w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8390w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8504w8754w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8504w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8510w8762w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8510w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8516w8770w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8516w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8521w8778w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8521w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8334w8786w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8334w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8340w8794w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8340w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8342w8802w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8342w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8344w8810w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8344w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8346w8818w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8346w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8348w8826w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8348w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8396w8610w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8396w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8350w8834w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8350w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8352w8842w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8352w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8354w8850w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8354w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8356w8858w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8356w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8402w8618w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8402w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8408w8626w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8408w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8414w8634w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8414w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8420w8642w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8420w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8426w8650w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8426w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8432w8658w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8432w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8438w8666w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8438w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9196w9394w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9196w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9255w9476w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9255w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9261w9484w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9261w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9267w9492w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9267w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9273w9500w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9273w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9279w9508w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9279w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9285w9516w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9285w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9291w9524w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9291w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9297w9532w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9297w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9303w9540w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9303w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9309w9548w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9309w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9201w9404w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9201w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9315w9556w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9315w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9321w9564w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9321w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9326w9572w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9326w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9141w9580w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9141w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9147w9588w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9147w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9149w9596w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9149w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9151w9604w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9151w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9153w9612w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9153w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9155w9620w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9155w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9157w9628w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9157w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9207w9412w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9207w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9159w9636w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9159w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9161w9644w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9161w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9163w9652w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9163w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9165w9660w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9165w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9213w9420w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9213w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9219w9428w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9219w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9225w9436w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9225w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9231w9444w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9231w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9237w9452w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9237w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9243w9460w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9243w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9249w9468w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9249w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10002w10191w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10002w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10061w10273w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10061w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10067w10281w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10067w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10073w10289w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10073w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10079w10297w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10079w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10085w10305w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10085w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10091w10313w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10091w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10097w10321w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10097w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10103w10329w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10103w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10109w10337w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10109w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10115w10345w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10115w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10007w10201w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10007w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10121w10353w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10121w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10126w10361w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10126w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9943w10369w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9943w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9949w10377w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9949w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9951w10385w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9951w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9953w10393w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9953w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9955w10401w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9955w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9957w10409w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9957w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9959w10417w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9959w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9961w10425w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9961w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10013w10209w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10013w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9963w10433w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9963w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9965w10441w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9965w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9967w10449w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9967w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9969w10457w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9969w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10019w10217w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10019w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10025w10225w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10025w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10031w10233w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10031w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10037w10241w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10037w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10043w10249w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10043w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10049w10257w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10049w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10055w10265w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10055w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range861w1149w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range861w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range920w1231w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range920w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range926w1239w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range926w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range932w1247w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range932w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range938w1255w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range938w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range944w1263w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range944w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range950w1271w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range950w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range956w1279w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range956w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range962w1287w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range962w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range968w1295w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range968w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range974w1303w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range974w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range866w1159w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range866w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range980w1311w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range980w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range986w1319w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range986w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range992w1327w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range992w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range998w1335w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range998w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1004w1343w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range1004w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1010w1351w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range1010w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1016w1359w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range1016w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1022w1367w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range1022w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1028w1375w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range1028w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1034w1383w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range1034w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range872w1167w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range872w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1040w1391w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range1040w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1046w1399w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range1046w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1051w1407w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range1051w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range846w1415w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range846w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range878w1175w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range878w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range884w1183w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range884w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range890w1191w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range890w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range896w1199w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range896w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range902w1207w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range902w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range908w1215w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range908w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range914w1223w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range914w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1717w1996w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1717w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1776w2078w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1776w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1782w2086w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1782w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1788w2094w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1788w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1794w2102w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1794w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1800w2110w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1800w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1806w2118w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1806w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1812w2126w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1812w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1818w2134w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1818w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1824w2142w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1824w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1830w2150w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1830w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1722w2006w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1722w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1836w2158w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1836w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1842w2166w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1842w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1848w2174w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1848w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1854w2182w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1854w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1860w2190w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1860w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1866w2198w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1866w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1872w2206w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1872w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1878w2214w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1878w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1884w2222w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1884w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1890w2230w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1890w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1728w2014w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1728w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1896w2238w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1896w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1901w2246w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1901w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1698w2254w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1698w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1704w2262w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1704w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1734w2022w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1734w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1740w2030w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1740w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1746w2038w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1746w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1752w2046w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1752w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1758w2054w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1758w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1764w2062w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1764w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1770w2070w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1770w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2568w2838w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2568w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2627w2920w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2627w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2633w2928w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2633w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2639w2936w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2639w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2645w2944w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2645w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2651w2952w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2651w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2657w2960w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2657w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2663w2968w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2663w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2669w2976w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2669w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2675w2984w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2675w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2681w2992w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2681w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2573w2848w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2573w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2687w3000w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2687w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2693w3008w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2693w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2699w3016w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2699w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2705w3024w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2705w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2711w3032w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2711w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2717w3040w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2717w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2723w3048w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2723w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2729w3056w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2729w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2735w3064w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2735w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2741w3072w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2741w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2579w2856w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2579w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2746w3080w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2746w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2545w3088w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2545w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2551w3096w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2551w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2553w3104w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2553w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2585w2864w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2585w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2591w2872w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2591w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2597w2880w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2597w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2603w2888w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2603w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2609w2896w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2609w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2615w2904w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2615w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2621w2912w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2621w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3414w3675w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3414w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3473w3757w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3473w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3479w3765w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3479w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3485w3773w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3485w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3491w3781w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3491w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3497w3789w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3497w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3503w3797w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3503w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3509w3805w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3509w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3515w3813w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3515w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3521w3821w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3521w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3527w3829w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3527w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3419w3685w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3419w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3533w3837w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3533w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3539w3845w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3539w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3545w3853w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3545w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3551w3861w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3551w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3557w3869w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3557w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3563w3877w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3563w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3569w3885w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3569w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3575w3893w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3575w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3581w3901w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3581w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3586w3909w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3586w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3425w3693w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3425w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3387w3917w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3387w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3393w3925w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3393w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3395w3933w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3395w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3397w3941w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3397w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3431w3701w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3431w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3437w3709w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3437w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3443w3717w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3443w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3449w3725w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3449w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3455w3733w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3455w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3461w3741w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3461w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3467w3749w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3467w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4255w4507w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4255w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4314w4589w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4314w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4320w4597w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4320w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4326w4605w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4326w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4332w4613w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4332w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4338w4621w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4338w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4344w4629w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4344w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4350w4637w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4350w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4356w4645w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4356w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4362w4653w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4362w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4368w4661w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4368w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4260w4517w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4260w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4374w4669w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4374w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4380w4677w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4380w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4386w4685w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4386w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4392w4693w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4392w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4398w4701w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4398w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4404w4709w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4404w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4410w4717w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4410w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4416w4725w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4416w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4421w4733w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4421w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4224w4741w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4224w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4266w4525w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4266w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4230w4749w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4230w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4232w4757w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4232w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4234w4765w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4234w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4236w4773w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4236w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4272w4533w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4272w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4278w4541w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4278w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4284w4549w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4284w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4290w4557w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4290w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4296w4565w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4296w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4302w4573w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4302w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4308w4581w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4308w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5091w5334w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5091w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5150w5416w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5150w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5156w5424w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5156w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5162w5432w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5162w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5168w5440w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5168w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5174w5448w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5174w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5180w5456w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5180w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5186w5464w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5186w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5192w5472w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5192w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5198w5480w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5198w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5204w5488w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5204w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5096w5344w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5096w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5210w5496w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5210w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5216w5504w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5216w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5222w5512w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5222w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5228w5520w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5228w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5234w5528w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5234w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5240w5536w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5240w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5246w5544w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5246w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5251w5552w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5251w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5056w5560w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5056w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5062w5568w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5062w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5102w5352w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5102w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5064w5576w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5064w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5066w5584w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5066w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5068w5592w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5068w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5070w5600w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5070w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5108w5360w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5108w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5114w5368w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5114w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5120w5376w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5120w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5126w5384w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5126w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5132w5392w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5132w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5138w5400w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5138w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5144w5408w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5144w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5922w6156w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5922w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5981w6238w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5981w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5987w6246w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5987w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5993w6254w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5993w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5999w6262w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5999w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6005w6270w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6005w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6011w6278w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6011w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6017w6286w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6017w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6023w6294w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6023w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6029w6302w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6029w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6035w6310w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6035w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5927w6166w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5927w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6041w6318w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6041w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6047w6326w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6047w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6053w6334w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6053w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6059w6342w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6059w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6065w6350w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6065w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6071w6358w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6071w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6076w6366w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6076w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5883w6374w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5883w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5889w6382w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5889w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5891w6390w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5891w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5933w6174w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5933w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5893w6398w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5893w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5895w6406w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5895w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5897w6414w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5897w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5899w6422w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5899w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5939w6182w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5939w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5945w6190w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5945w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5951w6198w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5951w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5957w6206w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5957w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5963w6214w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5963w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5969w6222w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5969w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5975w6230w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5975w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6748w6973w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6748w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6807w7055w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6807w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6813w7063w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6813w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6819w7071w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6819w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6825w7079w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6825w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6831w7087w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6831w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6837w7095w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6837w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6843w7103w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6843w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6849w7111w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6849w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6855w7119w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6855w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6861w7127w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6861w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6753w6983w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6753w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6867w7135w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6867w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6873w7143w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6873w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6879w7151w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6879w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6885w7159w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6885w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6891w7167w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6891w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6896w7175w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6896w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6705w7183w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6705w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6711w7191w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6711w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6713w7199w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6713w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6715w7207w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6715w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6759w6991w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6759w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6717w7215w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6717w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6719w7223w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6719w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6721w7231w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6721w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6723w7239w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6723w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6765w6999w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6765w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6771w7007w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6771w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6777w7015w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6777w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6783w7023w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6783w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6789w7031w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6789w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6795w7039w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6795w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6801w7047w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6801w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7714w7783w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7714w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7743w7866w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7743w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7746w7874w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7746w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7749w7882w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7749w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7752w7890w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7752w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7755w7898w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7755w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7758w7906w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7758w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7761w7914w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7761w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7764w7922w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7764w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7767w7930w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7767w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7770w7938w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7770w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7716w7794w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7716w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7773w7946w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7773w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7776w7954w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7776w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7779w7962w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7779w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7544w7970w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7544w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7548w7978w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7548w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7550w7986w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7550w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7552w7994w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7552w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7554w8002w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7554w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7556w8010w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7556w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7558w8018w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7558w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7719w7802w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7719w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7560w8026w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7560w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7562w8034w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7562w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7564w8042w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7564w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7566w8050w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7566w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7722w7810w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7722w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7725w7818w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7725w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7728w7826w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7728w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7731w7834w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7731w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7734w7842w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7734w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7737w7850w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7737w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7740w7858w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7740w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8524w8590w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8524w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8553w8673w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8553w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8556w8681w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8556w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8559w8689w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8559w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8562w8697w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8562w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8565w8705w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8565w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8568w8713w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8568w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8571w8721w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8571w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8574w8729w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8574w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8577w8737w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8577w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8580w8745w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8580w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8526w8601w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8526w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8583w8753w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8583w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8586w8761w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8586w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8358w8769w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8358w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8362w8777w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8362w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8364w8785w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8364w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8366w8793w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8366w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8368w8801w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8368w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8370w8809w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8370w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8372w8817w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8372w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8374w8825w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8374w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8529w8609w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8529w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8376w8833w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8376w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8378w8841w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8378w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8380w8849w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8380w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8382w8857w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8382w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8532w8617w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8532w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8535w8625w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8535w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8538w8633w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8538w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8541w8641w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8541w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8544w8649w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8544w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8547w8657w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8547w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8550w8665w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8550w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9329w9392w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9329w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9358w9475w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9358w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9361w9483w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9361w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9364w9491w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9364w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9367w9499w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9367w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9370w9507w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9370w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9373w9515w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9373w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9376w9523w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9376w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9379w9531w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9379w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9382w9539w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9382w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9385w9547w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9385w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9331w9403w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9331w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9388w9555w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9388w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9167w9563w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9167w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9171w9571w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9171w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9173w9579w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9173w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9175w9587w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9175w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9177w9595w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9177w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9179w9603w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9179w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9181w9611w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9181w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9183w9619w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9183w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9185w9627w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9185w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9334w9411w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9334w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9187w9635w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9187w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9189w9643w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9189w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9191w9651w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9191w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9193w9659w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9193w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9337w9419w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9337w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9340w9427w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9340w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9343w9435w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9343w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9346w9443w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9346w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9349w9451w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9349w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9352w9459w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9352w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9355w9467w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9355w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10129w10189w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10129w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10158w10272w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10158w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10161w10280w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10161w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10164w10288w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10164w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10167w10296w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10167w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10170w10304w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10170w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10173w10312w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10173w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10176w10320w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10176w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10179w10328w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10179w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10182w10336w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10182w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10185w10344w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10185w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10131w10200w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10131w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9971w10352w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9971w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9975w10360w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9975w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9977w10368w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9977w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9979w10376w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9979w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9981w10384w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9981w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9983w10392w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9983w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9985w10400w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9985w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9987w10408w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9987w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9989w10416w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9989w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9991w10424w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9991w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10134w10208w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10134w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9993w10432w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9993w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9995w10440w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9995w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9997w10448w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9997w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9999w10456w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9999w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10137w10216w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10137w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10140w10224w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10140w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10143w10232w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10143w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10146w10240w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10146w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10149w10248w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10149w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10152w10256w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10152w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10155w10264w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10155w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1054w1147w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1054w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1083w1230w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1083w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1086w1238w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1086w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1089w1246w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1089w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1092w1254w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1092w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1095w1262w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1095w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1098w1270w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1098w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1101w1278w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1101w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1104w1286w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1104w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1107w1294w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1107w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1110w1302w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1110w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1056w1158w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1056w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1113w1310w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1113w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1116w1318w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1116w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1119w1326w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1119w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1122w1334w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1122w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1125w1342w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1125w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1128w1350w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1128w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1131w1358w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1131w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1134w1366w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1134w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1137w1374w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1137w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1140w1382w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1140w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1059w1166w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1059w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1143w1390w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1143w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range852w1398w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range852w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range856w1406w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range856w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range858w1414w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range858w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1062w1174w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1062w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1065w1182w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1065w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1068w1190w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1068w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1071w1198w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1071w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1074w1206w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1074w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1077w1214w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1077w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1080w1222w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1080w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1904w1994w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1904w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1933w2077w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1933w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1936w2085w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1936w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1939w2093w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1939w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1942w2101w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1942w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1945w2109w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1945w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1948w2117w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1948w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1951w2125w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1951w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1954w2133w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1954w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1957w2141w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1957w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1960w2149w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1960w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1906w2005w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1906w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1963w2157w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1963w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1966w2165w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1966w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1969w2173w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1969w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1972w2181w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1972w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1975w2189w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1975w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1978w2197w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1978w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1981w2205w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1981w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1984w2213w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1984w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1987w2221w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1987w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1990w2229w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1990w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1909w2013w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1909w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1706w2237w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1706w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1710w2245w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1710w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1712w2253w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1712w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1714w2261w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1714w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1912w2021w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1912w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1915w2029w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1915w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1918w2037w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1918w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1921w2045w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1921w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1924w2053w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1924w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1927w2061w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1927w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1930w2069w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1930w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2749w2836w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2749w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2778w2919w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2778w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2781w2927w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2781w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2784w2935w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2784w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2787w2943w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2787w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2790w2951w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2790w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2793w2959w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2793w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2796w2967w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2796w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2799w2975w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2799w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2802w2983w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2802w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2805w2991w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2805w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2751w2847w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2751w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2808w2999w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2808w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2811w3007w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2811w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2814w3015w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2814w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2817w3023w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2817w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2820w3031w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2820w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2823w3039w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2823w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2826w3047w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2826w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2829w3055w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2829w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2832w3063w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2832w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2555w3071w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2555w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2754w2855w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2754w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2559w3079w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2559w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2561w3087w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2561w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2563w3095w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2563w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2565w3103w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2565w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2757w2863w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2757w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2760w2871w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2760w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2763w2879w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2763w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2766w2887w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2766w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2769w2895w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2769w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2772w2903w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2772w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2775w2911w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2775w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3589w3673w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3589w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3618w3756w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3618w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3621w3764w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3621w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3624w3772w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3624w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3627w3780w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3627w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3630w3788w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3630w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3633w3796w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3633w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3636w3804w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3636w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3639w3812w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3639w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3642w3820w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3642w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3645w3828w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3645w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3591w3684w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3591w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3648w3836w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3648w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3651w3844w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3651w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3654w3852w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3654w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3657w3860w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3657w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3660w3868w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3660w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3663w3876w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3663w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3666w3884w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3666w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3669w3892w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3669w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3399w3900w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3399w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3403w3908w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3403w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3594w3692w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3594w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3405w3916w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3405w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3407w3924w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3407w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3409w3932w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3409w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3411w3940w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3411w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3597w3700w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3597w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3600w3708w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3600w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3603w3716w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3603w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3606w3724w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3606w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3609w3732w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3609w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3612w3740w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3612w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3615w3748w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3615w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4424w4505w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4424w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4453w4588w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4453w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4456w4596w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4456w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4459w4604w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4459w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4462w4612w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4462w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4465w4620w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4465w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4468w4628w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4468w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4471w4636w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4471w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4474w4644w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4474w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4477w4652w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4477w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4480w4660w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4480w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4426w4516w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4426w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4483w4668w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4483w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4486w4676w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4486w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4489w4684w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4489w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4492w4692w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4492w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4495w4700w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4495w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4498w4708w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4498w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4501w4716w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4501w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4238w4724w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4238w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4242w4732w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4242w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4244w4740w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4244w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4429w4524w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4429w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4246w4748w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4246w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4248w4756w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4248w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4250w4764w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4250w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4252w4772w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4252w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4432w4532w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4432w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4435w4540w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4435w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4438w4548w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4438w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4441w4556w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4441w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4444w4564w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4444w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4447w4572w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4447w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4450w4580w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4450w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5254w5332w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5254w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5283w5415w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5283w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5286w5423w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5286w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5289w5431w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5289w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5292w5439w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5292w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5295w5447w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5295w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5298w5455w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5298w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5301w5463w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5301w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5304w5471w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5304w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5307w5479w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5307w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5310w5487w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5310w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5256w5343w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5256w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5313w5495w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5313w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5316w5503w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5316w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5319w5511w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5319w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5322w5519w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5322w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5325w5527w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5325w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5328w5535w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5328w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5072w5543w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5072w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5076w5551w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5076w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5078w5559w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5078w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5080w5567w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5080w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5259w5351w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5259w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5082w5575w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5082w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5084w5583w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5084w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5086w5591w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5086w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5088w5599w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5088w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5262w5359w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5262w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5265w5367w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5265w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5268w5375w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5268w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5271w5383w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5271w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5274w5391w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5274w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5277w5399w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5277w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5280w5407w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5280w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6079w6154w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6079w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6108w6237w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6108w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6111w6245w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6111w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6114w6253w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6114w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6117w6261w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6117w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6120w6269w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6120w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6123w6277w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6123w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6126w6285w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6126w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6129w6293w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6129w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6132w6301w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6132w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6135w6309w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6135w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6081w6165w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6081w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6138w6317w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6138w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6141w6325w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6141w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6144w6333w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6144w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6147w6341w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6147w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6150w6349w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6150w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5901w6357w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5901w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5905w6365w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5905w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5907w6373w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5907w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5909w6381w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5909w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5911w6389w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5911w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6084w6173w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6084w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5913w6397w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5913w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5915w6405w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5915w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5917w6413w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5917w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5919w6421w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5919w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6087w6181w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6087w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6090w6189w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6090w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6093w6197w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6093w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6096w6205w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6096w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6099w6213w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6099w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6102w6221w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6102w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6105w6229w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6105w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6899w6971w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6899w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6928w7054w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6928w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6931w7062w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6931w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6934w7070w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6934w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6937w7078w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6937w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6940w7086w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6940w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6943w7094w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6943w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6946w7102w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6946w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6949w7110w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6949w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6952w7118w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6952w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6955w7126w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6955w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6901w6982w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6901w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6958w7134w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6958w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6961w7142w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6961w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6964w7150w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6964w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6967w7158w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6967w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6725w7166w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6725w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6729w7174w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6729w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6731w7182w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6731w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6733w7190w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6733w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6735w7198w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6735w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6737w7206w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6737w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6904w6990w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6904w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6739w7214w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6739w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6741w7222w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6741w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6743w7230w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6743w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6745w7238w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6745w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6907w6998w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6907w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6910w7006w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6910w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6913w7014w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6913w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6916w7022w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6916w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6919w7030w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6919w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6922w7038w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6922w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6925w7046w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6925w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7572w7790w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7572w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7631w7871w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7631w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7637w7879w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7637w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7643w7887w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7643w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7649w7895w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7649w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7655w7903w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7655w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7661w7911w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7661w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7667w7919w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7667w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7673w7927w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7673w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7679w7935w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7679w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7685w7943w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7685w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7577w7799w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7577w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7691w7951w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7691w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7697w7959w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7697w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7703w7967w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7703w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7709w7975w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7709w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7712w7983w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7712w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7526w7991w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7526w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7529w7999w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7529w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7531w8007w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7531w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7533w8015w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7533w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7535w8023w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7535w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7583w7807w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7583w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7537w8031w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7537w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7539w8039w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7539w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7541w8047w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7541w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7543w8055w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7543w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7589w7815w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7589w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7595w7823w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7595w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7601w7831w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7601w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7607w7839w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7607w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7613w7847w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7613w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7619w7855w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7619w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7625w7863w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7625w(0) AND wire_indexbitff_w_lg_w_q_range607w7784w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8388w8597w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8388w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8447w8678w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8447w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8453w8686w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8453w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8459w8694w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8459w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8465w8702w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8465w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8471w8710w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8471w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8477w8718w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8477w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8483w8726w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8483w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8489w8734w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8489w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8495w8742w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8495w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8501w8750w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8501w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8393w8606w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8393w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8507w8758w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8507w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8513w8766w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8513w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8519w8774w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8519w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8522w8782w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8522w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8338w8790w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8338w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8341w8798w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8341w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8343w8806w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8343w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8345w8814w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8345w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8347w8822w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8347w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8349w8830w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8349w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8399w8614w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8399w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8351w8838w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8351w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8353w8846w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8353w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8355w8854w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8355w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8357w8862w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8357w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8405w8622w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8405w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8411w8630w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8411w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8417w8638w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8417w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8423w8646w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8423w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8429w8654w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8429w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8435w8662w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8435w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8441w8670w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8441w(0) AND wire_indexbitff_w_lg_w_q_range610w8591w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9199w9399w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9199w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9258w9480w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9258w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9264w9488w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9264w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9270w9496w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9270w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9276w9504w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9276w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9282w9512w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9282w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9288w9520w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9288w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9294w9528w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9294w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9300w9536w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9300w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9306w9544w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9306w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9312w9552w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9312w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9204w9408w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9204w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9318w9560w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9318w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9324w9568w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9324w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9327w9576w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9327w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9145w9584w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9145w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9148w9592w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9148w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9150w9600w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9150w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9152w9608w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9152w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9154w9616w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9154w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9156w9624w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9156w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9158w9632w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9158w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9210w9416w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9210w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9160w9640w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9160w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9162w9648w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9162w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9164w9656w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9164w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9166w9664w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9166w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9216w9424w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9216w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9222w9432w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9222w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9228w9440w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9228w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9234w9448w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9234w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9240w9456w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9240w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9246w9464w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9246w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9252w9472w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9252w(0) AND wire_indexbitff_w_lg_w_q_range613w9393w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10005w10196w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10005w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10064w10277w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10064w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10070w10285w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10070w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10076w10293w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10076w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10082w10301w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10082w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10088w10309w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10088w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10094w10317w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10094w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10100w10325w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10100w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10106w10333w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10106w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10112w10341w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10112w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10118w10349w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10118w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10010w10205w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10010w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10124w10357w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10124w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10127w10365w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10127w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9947w10373w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9947w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9950w10381w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9950w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9952w10389w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9952w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9954w10397w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9954w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9956w10405w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9956w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9958w10413w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9958w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9960w10421w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9960w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9962w10429w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9962w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10016w10213w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10016w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9964w10437w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9964w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9966w10445w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9966w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9968w10453w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9968w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9970w10461w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9970w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10022w10221w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10022w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10028w10229w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10028w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10034w10237w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10034w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10040w10245w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10040w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10046w10253w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10046w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10052w10261w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10052w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10058w10269w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10058w(0) AND wire_indexbitff_w_lg_w_q_range616w10190w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range864w1154w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range864w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range923w1235w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range923w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range929w1243w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range929w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range935w1251w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range935w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range941w1259w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range941w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range947w1267w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range947w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range953w1275w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range953w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range959w1283w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range959w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range965w1291w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range965w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range971w1299w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range971w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range977w1307w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range977w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range869w1163w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range869w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range983w1315w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range983w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range989w1323w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range989w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range995w1331w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range995w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1001w1339w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range1001w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1007w1347w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range1007w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1013w1355w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range1013w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1019w1363w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range1019w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1025w1371w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range1025w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1031w1379w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range1031w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1037w1387w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range1037w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range875w1171w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range875w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1043w1395w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range1043w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1049w1403w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range1049w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1052w1411w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range1052w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range850w1419w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range850w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range881w1179w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range881w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range887w1187w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range887w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range893w1195w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range893w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range899w1203w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range899w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range905w1211w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range905w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range911w1219w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range911w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range917w1227w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range917w(0) AND wire_indexbitff_w_lg_w_q_range583w1148w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1720w2001w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1720w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1779w2082w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1779w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1785w2090w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1785w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1791w2098w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1791w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1797w2106w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1797w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1803w2114w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1803w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1809w2122w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1809w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1815w2130w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1815w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1821w2138w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1821w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1827w2146w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1827w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1833w2154w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1833w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1725w2010w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1725w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1839w2162w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1839w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1845w2170w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1845w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1851w2178w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1851w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1857w2186w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1857w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1863w2194w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1863w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1869w2202w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1869w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1875w2210w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1875w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1881w2218w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1881w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1887w2226w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1887w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1893w2234w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1893w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1731w2018w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1731w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1899w2242w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1899w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1902w2250w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1902w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1702w2258w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1702w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1705w2266w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1705w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1737w2026w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1737w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1743w2034w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1743w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1749w2042w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1749w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1755w2050w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1755w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1761w2058w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1761w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1767w2066w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1767w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1773w2074w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1773w(0) AND wire_indexbitff_w_lg_w_q_range586w1995w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2571w2843w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2571w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2630w2924w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2630w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2636w2932w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2636w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2642w2940w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2642w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2648w2948w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2648w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2654w2956w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2654w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2660w2964w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2660w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2666w2972w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2666w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2672w2980w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2672w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2678w2988w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2678w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2684w2996w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2684w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2576w2852w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2576w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2690w3004w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2690w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2696w3012w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2696w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2702w3020w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2702w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2708w3028w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2708w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2714w3036w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2714w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2720w3044w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2720w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2726w3052w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2726w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2732w3060w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2732w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2738w3068w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2738w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2744w3076w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2744w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2582w2860w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2582w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2747w3084w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2747w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2549w3092w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2549w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2552w3100w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2552w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2554w3108w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2554w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2588w2868w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2588w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2594w2876w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2594w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2600w2884w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2600w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2606w2892w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2606w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2612w2900w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2612w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2618w2908w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2618w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2624w2916w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2624w(0) AND wire_indexbitff_w_lg_w_q_range589w2837w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3417w3680w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3417w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3476w3761w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3476w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3482w3769w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3482w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3488w3777w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3488w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3494w3785w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3494w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3500w3793w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3500w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3506w3801w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3506w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3512w3809w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3512w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3518w3817w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3518w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3524w3825w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3524w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3530w3833w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3530w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3422w3689w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3422w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3536w3841w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3536w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3542w3849w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3542w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3548w3857w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3548w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3554w3865w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3554w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3560w3873w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3560w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3566w3881w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3566w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3572w3889w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3572w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3578w3897w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3578w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3584w3905w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3584w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3587w3913w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3587w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3428w3697w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3428w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3391w3921w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3391w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3394w3929w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3394w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3396w3937w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3396w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3398w3945w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3398w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3434w3705w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3434w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3440w3713w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3440w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3446w3721w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3446w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3452w3729w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3452w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3458w3737w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3458w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3464w3745w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3464w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3470w3753w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3470w(0) AND wire_indexbitff_w_lg_w_q_range592w3674w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4258w4512w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4258w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4317w4593w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4317w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4323w4601w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4323w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4329w4609w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4329w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4335w4617w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4335w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4341w4625w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4341w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4347w4633w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4347w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4353w4641w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4353w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4359w4649w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4359w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4365w4657w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4365w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4371w4665w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4371w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4263w4521w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4263w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4377w4673w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4377w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4383w4681w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4383w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4389w4689w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4389w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4395w4697w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4395w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4401w4705w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4401w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4407w4713w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4407w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4413w4721w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4413w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4419w4729w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4419w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4422w4737w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4422w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4228w4745w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4228w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4269w4529w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4269w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4231w4753w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4231w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4233w4761w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4233w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4235w4769w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4235w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4237w4777w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4237w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4275w4537w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4275w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4281w4545w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4281w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4287w4553w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4287w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4293w4561w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4293w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4299w4569w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4299w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4305w4577w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4305w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4311w4585w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4311w(0) AND wire_indexbitff_w_lg_w_q_range595w4506w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5094w5339w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5094w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5153w5420w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5153w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5159w5428w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5159w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5165w5436w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5165w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5171w5444w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5171w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5177w5452w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5177w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5183w5460w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5183w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5189w5468w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5189w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5195w5476w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5195w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5201w5484w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5201w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5207w5492w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5207w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5099w5348w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5099w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5213w5500w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5213w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5219w5508w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5219w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5225w5516w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5225w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5231w5524w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5231w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5237w5532w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5237w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5243w5540w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5243w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5249w5548w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5249w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5252w5556w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5252w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5060w5564w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5060w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5063w5572w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5063w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5105w5356w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5105w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5065w5580w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5065w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5067w5588w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5067w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5069w5596w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5069w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5071w5604w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5071w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5111w5364w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5111w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5117w5372w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5117w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5123w5380w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5123w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5129w5388w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5129w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5135w5396w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5135w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5141w5404w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5141w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5147w5412w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5147w(0) AND wire_indexbitff_w_lg_w_q_range598w5333w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5925w6161w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5925w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5984w6242w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5984w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5990w6250w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5990w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5996w6258w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5996w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6002w6266w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6002w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6008w6274w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6008w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6014w6282w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6014w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6020w6290w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6020w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6026w6298w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6026w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6032w6306w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6032w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6038w6314w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6038w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5930w6170w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5930w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6044w6322w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6044w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6050w6330w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6050w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6056w6338w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6056w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6062w6346w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6062w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6068w6354w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6068w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6074w6362w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6074w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6077w6370w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6077w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5887w6378w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5887w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5890w6386w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5890w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5892w6394w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5892w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5936w6178w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5936w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5894w6402w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5894w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5896w6410w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5896w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5898w6418w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5898w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5900w6426w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5900w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5942w6186w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5942w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5948w6194w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5948w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5954w6202w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5954w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5960w6210w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5960w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5966w6218w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5966w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5972w6226w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5972w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5978w6234w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5978w(0) AND wire_indexbitff_w_lg_w_q_range601w6155w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6751w6978w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6751w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6810w7059w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6810w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6816w7067w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6816w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6822w7075w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6822w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6828w7083w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6828w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6834w7091w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6834w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6840w7099w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6840w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6846w7107w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6846w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6852w7115w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6852w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6858w7123w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6858w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6864w7131w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6864w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6756w6987w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6756w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6870w7139w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6870w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6876w7147w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6876w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6882w7155w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6882w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6888w7163w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6888w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6894w7171w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6894w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6897w7179w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6897w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6709w7187w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6709w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6712w7195w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6712w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6714w7203w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6714w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6716w7211w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6716w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6762w6995w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6762w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6718w7219w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6718w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6720w7227w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6720w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6722w7235w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6722w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6724w7243w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6724w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6768w7003w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6768w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6774w7011w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6774w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6780w7019w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6780w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6786w7027w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6786w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6792w7035w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6792w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6798w7043w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6798w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6804w7051w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6804w(0) AND wire_indexbitff_w_lg_w_q_range604w6972w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7715w7789w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7715w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7744w7870w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7744w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7747w7878w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7747w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7750w7886w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7750w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7753w7894w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7753w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7756w7902w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7756w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7759w7910w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7759w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7762w7918w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7762w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7765w7926w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7765w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7768w7934w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7768w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7771w7942w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7771w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7717w7798w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7717w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7774w7950w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7774w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7777w7958w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7777w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7780w7966w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7780w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7546w7974w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7546w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7549w7982w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7549w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7551w7990w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7551w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7553w7998w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7553w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7555w8006w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7555w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7557w8014w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7557w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7559w8022w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7559w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7720w7806w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7720w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7561w8030w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7561w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7563w8038w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7563w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7565w8046w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7565w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7567w8054w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7567w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7723w7814w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7723w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7726w7822w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7726w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7729w7830w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7729w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7732w7838w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7732w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7735w7846w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7735w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7738w7854w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7738w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7741w7862w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7741w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8525w8596w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8525w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8554w8677w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8554w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8557w8685w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8557w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8560w8693w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8560w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8563w8701w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8563w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8566w8709w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8566w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8569w8717w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8569w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8572w8725w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8572w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8575w8733w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8575w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8578w8741w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8578w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8581w8749w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8581w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8527w8605w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8527w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8584w8757w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8584w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8587w8765w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8587w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8360w8773w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8360w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8363w8781w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8363w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8365w8789w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8365w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8367w8797w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8367w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8369w8805w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8369w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8371w8813w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8371w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8373w8821w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8373w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8375w8829w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8375w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8530w8613w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8530w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8377w8837w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8377w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8379w8845w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8379w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8381w8853w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8381w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8383w8861w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8383w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8533w8621w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8533w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8536w8629w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8536w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8539w8637w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8539w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8542w8645w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8542w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8545w8653w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8545w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8548w8661w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8548w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8551w8669w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8551w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9330w9398w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9330w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9359w9479w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9359w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9362w9487w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9362w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9365w9495w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9365w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9368w9503w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9368w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9371w9511w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9371w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9374w9519w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9374w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9377w9527w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9377w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9380w9535w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9380w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9383w9543w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9383w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9386w9551w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9386w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9332w9407w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9332w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9389w9559w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9389w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9169w9567w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9169w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9172w9575w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9172w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9174w9583w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9174w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9176w9591w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9176w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9178w9599w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9178w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9180w9607w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9180w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9182w9615w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9182w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9184w9623w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9184w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9186w9631w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9186w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9335w9415w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9335w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9188w9639w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9188w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9190w9647w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9190w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9192w9655w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9192w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9194w9663w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9194w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9338w9423w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9338w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9341w9431w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9341w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9344w9439w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9344w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9347w9447w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9347w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9350w9455w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9350w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9353w9463w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9353w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9356w9471w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9356w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10130w10195w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10130w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10159w10276w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10159w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10162w10284w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10162w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10165w10292w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10165w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10168w10300w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10168w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10171w10308w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10171w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10174w10316w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10174w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10177w10324w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10177w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10180w10332w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10180w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10183w10340w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10183w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10186w10348w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10186w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10132w10204w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10132w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9973w10356w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9973w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9976w10364w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9976w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9978w10372w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9978w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9980w10380w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9980w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9982w10388w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9982w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9984w10396w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9984w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9986w10404w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9986w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9988w10412w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9988w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9990w10420w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9990w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9992w10428w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9992w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10135w10212w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10135w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9994w10436w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9994w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9996w10444w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9996w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9998w10452w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9998w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10000w10460w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10000w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10138w10220w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10138w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10141w10228w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10141w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10144w10236w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10144w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10147w10244w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10147w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10150w10252w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10150w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10153w10260w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10153w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10156w10268w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10156w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1055w1153w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1055w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1084w1234w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1084w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1087w1242w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1087w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1090w1250w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1090w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1093w1258w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1093w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1096w1266w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1096w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1099w1274w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1099w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1102w1282w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1102w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1105w1290w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1105w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1108w1298w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1108w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1111w1306w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1111w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1057w1162w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1057w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1114w1314w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1114w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1117w1322w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1117w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1120w1330w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1120w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1123w1338w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1123w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1126w1346w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1126w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1129w1354w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1129w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1132w1362w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1132w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1135w1370w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1135w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1138w1378w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1138w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1141w1386w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1141w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1060w1170w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1060w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1144w1394w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1144w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range854w1402w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range854w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range857w1410w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range857w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range859w1418w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range859w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1063w1178w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1063w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1066w1186w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1066w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1069w1194w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1069w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1072w1202w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1072w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1075w1210w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1075w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1078w1218w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1078w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1081w1226w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1081w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1905w2000w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1905w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1934w2081w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1934w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1937w2089w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1937w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1940w2097w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1940w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1943w2105w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1943w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1946w2113w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1946w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1949w2121w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1949w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1952w2129w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1952w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1955w2137w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1955w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1958w2145w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1958w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1961w2153w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1961w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1907w2009w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1907w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1964w2161w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1964w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1967w2169w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1967w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1970w2177w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1970w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1973w2185w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1973w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1976w2193w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1976w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1979w2201w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1979w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1982w2209w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1982w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1985w2217w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1985w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1988w2225w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1988w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1991w2233w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1991w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1910w2017w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1910w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1708w2241w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1708w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1711w2249w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1711w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1713w2257w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1713w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1715w2265w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1715w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1913w2025w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1913w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1916w2033w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1916w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1919w2041w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1919w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1922w2049w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1922w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1925w2057w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1925w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1928w2065w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1928w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1931w2073w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1931w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2750w2842w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2750w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2779w2923w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2779w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2782w2931w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2782w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2785w2939w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2785w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2788w2947w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2788w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2791w2955w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2791w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2794w2963w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2794w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2797w2971w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2797w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2800w2979w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2800w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2803w2987w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2803w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2806w2995w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2806w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2752w2851w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2752w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2809w3003w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2809w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2812w3011w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2812w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2815w3019w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2815w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2818w3027w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2818w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2821w3035w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2821w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2824w3043w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2824w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2827w3051w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2827w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2830w3059w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2830w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2833w3067w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2833w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2557w3075w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2557w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2755w2859w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2755w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2560w3083w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2560w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2562w3091w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2562w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2564w3099w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2564w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2566w3107w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2566w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2758w2867w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2758w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2761w2875w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2761w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2764w2883w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2764w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2767w2891w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2767w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2770w2899w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2770w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2773w2907w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2773w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2776w2915w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2776w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3590w3679w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3590w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3619w3760w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3619w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3622w3768w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3622w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3625w3776w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3625w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3628w3784w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3628w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3631w3792w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3631w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3634w3800w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3634w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3637w3808w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3637w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3640w3816w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3640w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3643w3824w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3643w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3646w3832w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3646w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3592w3688w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3592w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3649w3840w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3649w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3652w3848w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3652w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3655w3856w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3655w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3658w3864w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3658w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3661w3872w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3661w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3664w3880w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3664w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3667w3888w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3667w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3670w3896w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3670w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3401w3904w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3401w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3404w3912w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3404w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3595w3696w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3595w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3406w3920w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3406w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3408w3928w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3408w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3410w3936w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3410w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3412w3944w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3412w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3598w3704w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3598w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3601w3712w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3601w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3604w3720w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3604w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3607w3728w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3607w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3610w3736w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3610w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3613w3744w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3613w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3616w3752w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3616w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4425w4511w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4425w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4454w4592w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4454w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4457w4600w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4457w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4460w4608w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4460w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4463w4616w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4463w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4466w4624w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4466w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4469w4632w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4469w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4472w4640w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4472w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4475w4648w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4475w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4478w4656w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4478w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4481w4664w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4481w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4427w4520w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4427w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4484w4672w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4484w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4487w4680w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4487w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4490w4688w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4490w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4493w4696w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4493w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4496w4704w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4496w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4499w4712w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4499w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4502w4720w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4502w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4240w4728w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4240w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4243w4736w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4243w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4245w4744w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4245w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4430w4528w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4430w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4247w4752w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4247w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4249w4760w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4249w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4251w4768w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4251w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4253w4776w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4253w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4433w4536w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4433w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4436w4544w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4436w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4439w4552w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4439w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4442w4560w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4442w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4445w4568w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4445w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4448w4576w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4448w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4451w4584w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4451w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5255w5338w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5255w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5284w5419w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5284w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5287w5427w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5287w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5290w5435w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5290w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5293w5443w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5293w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5296w5451w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5296w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5299w5459w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5299w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5302w5467w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5302w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5305w5475w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5305w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5308w5483w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5308w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5311w5491w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5311w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5257w5347w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5257w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5314w5499w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5314w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5317w5507w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5317w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5320w5515w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5320w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5323w5523w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5323w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5326w5531w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5326w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5329w5539w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5329w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5074w5547w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5074w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5077w5555w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5077w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5079w5563w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5079w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5081w5571w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5081w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5260w5355w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5260w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5083w5579w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5083w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5085w5587w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5085w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5087w5595w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5087w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5089w5603w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5089w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5263w5363w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5263w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5266w5371w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5266w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5269w5379w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5269w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5272w5387w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5272w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5275w5395w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5275w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5278w5403w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5278w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5281w5411w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5281w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6080w6160w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6080w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6109w6241w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6109w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6112w6249w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6112w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6115w6257w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6115w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6118w6265w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6118w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6121w6273w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6121w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6124w6281w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6124w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6127w6289w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6127w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6130w6297w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6130w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6133w6305w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6133w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6136w6313w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6136w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6082w6169w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6082w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6139w6321w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6139w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6142w6329w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6142w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6145w6337w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6145w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6148w6345w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6148w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6151w6353w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6151w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5903w6361w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5903w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5906w6369w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5906w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5908w6377w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5908w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5910w6385w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5910w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5912w6393w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5912w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6085w6177w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6085w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5914w6401w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5914w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5916w6409w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5916w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5918w6417w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5918w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5920w6425w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5920w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6088w6185w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6088w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6091w6193w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6091w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6094w6201w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6094w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6097w6209w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6097w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6100w6217w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6100w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6103w6225w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6103w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6106w6233w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6106w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6900w6977w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6900w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6929w7058w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6929w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6932w7066w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6932w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6935w7074w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6935w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6938w7082w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6938w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6941w7090w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6941w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6944w7098w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6944w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6947w7106w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6947w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6950w7114w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6950w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6953w7122w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6953w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6956w7130w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6956w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6902w6986w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6902w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6959w7138w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6959w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6962w7146w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6962w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6965w7154w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6965w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6968w7162w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6968w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6727w7170w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6727w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6730w7178w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6730w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6732w7186w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6732w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6734w7194w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6734w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6736w7202w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6736w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6738w7210w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6738w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6905w6994w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6905w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6740w7218w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6740w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6742w7226w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6742w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6744w7234w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6744w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6746w7242w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6746w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6908w7002w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6908w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6911w7010w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6911w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6914w7018w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6914w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6917w7026w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6917w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6920w7034w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6920w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6923w7042w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6923w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6926w7050w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6926w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_indexbit412w(0) <= NOT indexbit;
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8871w8873w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8871w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8952w8954w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8952w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8960w8962w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8960w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8968w8970w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8968w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8976w8978w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8984w8986w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8984w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8992w8994w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8992w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9000w9002w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9000w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9008w9010w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9008w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9016w9018w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9016w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9024w9026w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9024w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8880w8882w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8880w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9032w9034w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9032w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9040w9042w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9040w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9048w9050w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9048w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9056w9058w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9056w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9064w9066w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9064w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9072w9074w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9072w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9080w9082w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9080w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9088w9090w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9088w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9096w9098w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9096w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9104w9106w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9104w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8888w8890w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8888w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9112w9114w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9112w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9120w9122w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9120w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9128w9130w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9128w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9136w9138w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9136w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8896w8898w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8896w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8904w8906w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8904w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8912w8914w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8912w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8920w8922w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8920w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8928w8930w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8928w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8936w8938w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8936w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8944w8946w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8944w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9673w9675w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9673w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9754w9756w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9754w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9762w9764w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9762w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9770w9772w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9770w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9778w9780w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9778w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9786w9788w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9786w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9794w9796w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9794w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9802w9804w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9802w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9810w9812w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9810w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9818w9820w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9818w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9826w9828w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9826w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9682w9684w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9682w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9834w9836w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9834w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9842w9844w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9842w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9850w9852w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9850w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9858w9860w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9858w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9866w9868w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9866w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9874w9876w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9874w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9882w9884w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9882w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9890w9892w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9890w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9898w9900w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9898w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9906w9908w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9906w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9690w9692w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9690w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9914w9916w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9914w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9922w9924w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9922w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9930w9932w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9930w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9938w9940w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9938w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9698w9700w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9698w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9706w9708w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9706w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9714w9716w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9714w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9722w9724w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9730w9732w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9730w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9738w9740w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9738w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9746w9748w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9746w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10470w10472w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10470w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10551w10553w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10551w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10559w10561w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10559w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10567w10569w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10567w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10575w10577w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10575w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10583w10585w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10583w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10591w10593w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10591w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10599w10601w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10599w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10607w10609w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10607w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10615w10617w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10615w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10623w10625w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10623w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10479w10481w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10479w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10631w10633w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10631w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10639w10641w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10639w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10647w10649w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10647w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10655w10657w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10655w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10663w10665w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10663w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10671w10673w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10671w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10679w10681w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10679w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10687w10689w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10687w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10695w10697w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10695w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10703w10705w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10703w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10487w10489w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10487w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10711w10713w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10711w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10719w10721w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10719w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10727w10729w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10727w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10735w10737w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10735w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10495w10497w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10495w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10503w10505w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10503w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10511w10513w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10511w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10519w10521w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10519w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10527w10529w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10527w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10535w10537w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10535w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10543w10545w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10543w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1428w1430w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1428w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1509w1511w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1509w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1517w1519w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1517w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1525w1527w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1525w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1533w1535w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1533w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1541w1543w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1541w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1549w1551w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1549w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1557w1559w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1557w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1565w1567w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1565w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1573w1575w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1573w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1581w1583w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1581w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1437w1439w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1437w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1589w1591w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1589w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1597w1599w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1597w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1605w1607w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1605w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1613w1615w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1613w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1621w1623w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1621w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1629w1631w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1629w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1637w1639w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1637w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1645w1647w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1645w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1653w1655w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1653w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1661w1663w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1661w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1445w1447w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1445w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1669w1671w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1669w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1677w1679w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1677w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1685w1687w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1685w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1693w1695w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1693w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1453w1455w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1453w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1461w1463w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1461w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1469w1471w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1469w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1477w1479w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1477w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1485w1487w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1485w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1493w1495w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1493w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1501w1503w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1501w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2275w2277w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2275w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2356w2358w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2356w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2364w2366w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2364w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2372w2374w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2372w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2380w2382w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2380w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2388w2390w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2388w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2396w2398w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2396w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2404w2406w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2404w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2412w2414w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2412w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2420w2422w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2420w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2428w2430w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2428w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2284w2286w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2284w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2436w2438w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2436w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2444w2446w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2444w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2452w2454w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2452w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2460w2462w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2460w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2468w2470w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2468w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2476w2478w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2476w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2484w2486w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2484w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2492w2494w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2492w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2500w2502w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2500w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2508w2510w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2508w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2292w2294w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2292w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2516w2518w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2516w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2524w2526w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2524w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2532w2534w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2532w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2540w2542w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2540w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2300w2302w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2300w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2308w2310w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2308w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2316w2318w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2316w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2324w2326w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2324w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2332w2334w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2332w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2340w2342w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2340w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2348w2350w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2348w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3117w3119w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3117w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3198w3200w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3198w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3206w3208w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3206w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3214w3216w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3214w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3222w3224w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3222w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3230w3232w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3230w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3238w3240w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3238w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3246w3248w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3246w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3254w3256w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3254w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3262w3264w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3262w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3270w3272w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3270w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3126w3128w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3126w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3278w3280w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3278w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3286w3288w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3286w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3294w3296w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3294w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3302w3304w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3302w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3310w3312w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3310w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3318w3320w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3318w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3326w3328w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3326w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3334w3336w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3334w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3342w3344w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3342w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3350w3352w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3350w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3134w3136w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3134w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3358w3360w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3358w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3366w3368w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3366w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3374w3376w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3374w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3382w3384w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3382w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3142w3144w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3142w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3150w3152w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3150w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3158w3160w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3158w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3166w3168w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3166w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3174w3176w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3174w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3182w3184w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3182w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3190w3192w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3190w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3954w3956w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3954w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4035w4037w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4035w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4043w4045w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4043w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4051w4053w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4051w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4059w4061w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4059w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4067w4069w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4067w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4075w4077w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4075w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4083w4085w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4083w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4091w4093w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4091w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4099w4101w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4099w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4107w4109w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4107w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3963w3965w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3963w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4115w4117w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4115w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4123w4125w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4123w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4131w4133w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4131w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4139w4141w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4139w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4147w4149w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4147w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4155w4157w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4155w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4163w4165w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4163w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4171w4173w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4171w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4179w4181w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4179w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4187w4189w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4187w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3971w3973w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3971w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4195w4197w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4195w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4203w4205w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4203w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4211w4213w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4211w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4219w4221w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4219w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3979w3981w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3979w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3987w3989w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3987w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3995w3997w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3995w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4003w4005w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4003w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4011w4013w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4011w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4019w4021w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4019w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4027w4029w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4027w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4786w4788w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4786w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4867w4869w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4867w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4875w4877w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4875w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4883w4885w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4883w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4891w4893w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4891w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4899w4901w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4899w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4907w4909w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4907w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4915w4917w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4915w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4923w4925w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4923w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4931w4933w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4931w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4939w4941w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4939w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4795w4797w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4795w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4947w4949w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4947w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4955w4957w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4955w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4963w4965w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4963w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4971w4973w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4971w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4979w4981w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4979w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4987w4989w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4987w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4995w4997w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4995w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5003w5005w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range5003w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5011w5013w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range5011w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5019w5021w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range5019w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4803w4805w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4803w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5027w5029w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range5027w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5035w5037w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range5035w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5043w5045w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range5043w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5051w5053w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range5051w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4811w4813w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4811w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4819w4821w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4819w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4827w4829w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4827w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4835w4837w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4835w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4843w4845w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4843w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4851w4853w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4851w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4859w4861w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4859w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5613w5615w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5613w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5694w5696w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5694w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5702w5704w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5702w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5710w5712w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5710w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5718w5720w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5718w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5726w5728w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5726w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5734w5736w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5734w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5742w5744w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5742w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5750w5752w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5750w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5758w5760w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5758w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5766w5768w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5766w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5622w5624w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5622w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5774w5776w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5774w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5782w5784w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5782w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5790w5792w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5790w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5798w5800w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5798w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5806w5808w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5806w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5814w5816w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5814w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5822w5824w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5822w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5830w5832w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5830w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5838w5840w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5838w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5846w5848w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5846w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5630w5632w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5630w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5854w5856w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5854w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5862w5864w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5862w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5870w5872w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5870w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5878w5880w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5878w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5638w5640w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5638w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5646w5648w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5646w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5654w5656w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5654w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5662w5664w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5662w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5670w5672w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5670w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5678w5680w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5678w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5686w5688w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5686w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6435w6437w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6435w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6516w6518w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6516w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6524w6526w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6524w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6532w6534w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6532w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6540w6542w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6540w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6548w6550w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6548w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6556w6558w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6556w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6564w6566w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6564w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6572w6574w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6572w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6580w6582w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6580w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6588w6590w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6588w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6444w6446w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6444w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6596w6598w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6596w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6604w6606w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6604w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6612w6614w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6612w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6620w6622w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6620w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6628w6630w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6628w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6636w6638w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6636w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6644w6646w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6644w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6652w6654w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6652w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6660w6662w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6660w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6668w6670w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6668w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6452w6454w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6452w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6676w6678w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6676w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6684w6686w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6684w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6692w6694w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6692w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6700w6702w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6700w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6460w6462w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6460w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6468w6470w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6468w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6476w6478w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6476w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6484w6486w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6484w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6492w6494w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6492w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6500w6502w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6500w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6508w6510w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6508w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7252w7254w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7252w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7333w7335w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7333w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7341w7343w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7341w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7349w7351w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7349w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7357w7359w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7357w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7365w7367w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7365w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7373w7375w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7373w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7381w7383w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7381w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7389w7391w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7389w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7397w7399w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7397w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7405w7407w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7405w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7261w7263w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7261w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7413w7415w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7413w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7421w7423w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7421w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7429w7431w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7429w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7437w7439w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7437w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7445w7447w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7445w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7453w7455w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7453w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7461w7463w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7461w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7469w7471w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7477w7479w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7477w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7485w7487w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7485w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7269w7271w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7269w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7493w7495w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7493w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7501w7503w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7501w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7509w7511w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7509w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7517w7519w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7517w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7277w7279w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7277w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7285w7287w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7285w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7293w7295w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7293w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7301w7303w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7301w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7309w7311w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7309w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7317w7319w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7317w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7325w7327w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7325w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8064w8066w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8064w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8145w8147w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8145w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8153w8155w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8153w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8161w8163w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8161w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8169w8171w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8169w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8177w8179w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8177w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8185w8187w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8185w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8193w8195w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8193w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8201w8203w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8201w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8209w8211w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8209w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8217w8219w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8217w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8073w8075w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8073w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8225w8227w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8233w8235w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8233w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8241w8243w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8241w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8249w8251w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8249w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8257w8259w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8257w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8265w8267w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8265w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8273w8275w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8273w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8281w8283w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8281w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8289w8291w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8289w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8297w8299w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8297w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8081w8083w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8081w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8305w8307w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8305w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8313w8315w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8313w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8321w8323w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8321w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8329w8331w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8329w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8089w8091w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8089w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8097w8099w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8097w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8105w8107w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8105w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8113w8115w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8113w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8121w8123w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8121w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8129w8131w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8129w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8137w8139w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8137w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10751w10755w10756w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10751w10755w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10750w10753w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10794w10807w10808w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10794w10807w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10804w10806w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10799w10812w10813w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10799w10812w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10809w10811w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10804w10817w10818w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10804w10817w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10814w10816w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10809w10822w10823w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10809w10822w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10819w10821w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10814w10827w10828w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10814w10827w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10824w10826w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10819w10832w10833w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10819w10832w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10829w10831w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10824w10837w10838w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10824w10837w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10834w10836w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10829w10842w10843w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10829w10842w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10839w10841w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10834w10847w10848w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10834w10847w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10844w10846w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10839w10852w10853w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10839w10852w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10849w10851w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10759w10762w10763w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10759w10762w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10758w10761w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10844w10857w10858w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10844w10857w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10854w10856w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10849w10862w10863w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10849w10862w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10859w10861w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10854w10867w10868w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10854w10867w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10864w10866w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10859w10872w10873w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10859w10872w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10869w10871w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10864w10877w10878w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10864w10877w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10874w10876w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10869w10882w10883w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10869w10882w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10879w10881w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10874w10887w10888w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10874w10887w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10884w10886w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10879w10892w10893w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10879w10892w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10889w10891w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10884w10897w10898w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10884w10897w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10894w10896w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10889w10902w10903w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10889w10902w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10899w10901w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10750w10767w10768w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10750w10767w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10764w10766w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10894w10907w10908w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10894w10907w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10904w10906w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10899w10912w10913w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10899w10912w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10909w10911w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10904w10915w10916w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10904w10915w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10909w10911w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10909w10918w10919w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10909w10918w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10909w10911w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10758w10772w10773w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10758w10772w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10769w10771w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10764w10777w10778w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10764w10777w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10774w10776w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10769w10782w10783w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10769w10782w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10779w10781w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10774w10787w10788w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10774w10787w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10784w10786w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10779w10792w10793w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10779w10792w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10789w10791w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10784w10797w10798w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10784w10797w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10794w10796w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10789w10802w10803w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10789w10802w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10799w10801w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range458w461w462w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range458w461w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range448w460w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range463w466w467w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range463w466w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range453w465w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range468w471w472w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range468w471w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range458w470w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range473w476w477w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range473w476w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range463w475w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range478w481w482w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range478w481w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range468w480w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range483w486w487w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range483w486w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range473w485w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range488w491w492w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range488w491w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range478w490w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range493w496w497w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range493w496w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range483w495w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range498w501w502w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range498w501w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range488w500w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range503w506w507w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range503w506w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range493w505w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range508w511w512w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range508w511w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range498w510w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range513w516w517w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range513w516w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range503w515w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range518w521w522w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range518w521w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range508w520w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range523w526w527w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range523w526w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range513w525w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range528w531w532w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range528w531w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range518w530w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range533w536w537w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range533w536w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range523w535w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range538w541w542w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range538w541w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range528w540w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range543w546w547w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range543w546w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range533w545w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range548w551w552w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range548w551w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range538w550w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range553w556w557w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range553w556w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range543w555w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range418w421w422w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range418w421w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range410w420w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range558w561w562w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range558w561w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range548w560w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range563w566w567w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range563w566w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range553w565w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range568w571w572w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range568w571w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range558w570w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range573w576w577w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range573w576w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range563w575w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range423w426w427w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range423w426w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range415w425w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range428w431w432w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range428w431w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range418w430w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range433w436w437w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range433w436w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range423w435w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range438w441w442w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range438w441w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range428w440w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range443w446w447w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range443w446w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range433w445w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range448w451w452w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range448w451w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range438w450w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range453w456w457w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range453w456w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range443w455w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7569w7785w7786w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7569w7785w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7714w7783w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7628w7867w7868w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7628w7867w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7743w7866w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7634w7875w7876w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7634w7875w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7746w7874w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7640w7883w7884w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7640w7883w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7749w7882w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7646w7891w7892w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7646w7891w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7752w7890w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7652w7899w7900w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7652w7899w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7755w7898w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7658w7907w7908w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7658w7907w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7758w7906w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7664w7915w7916w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7664w7915w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7761w7914w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7670w7923w7924w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7670w7923w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7764w7922w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7676w7931w7932w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7676w7931w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7767w7930w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7682w7939w7940w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7682w7939w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7770w7938w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7574w7795w7796w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7574w7795w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7716w7794w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7688w7947w7948w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7688w7947w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7773w7946w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7694w7955w7956w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7694w7955w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7776w7954w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7700w7963w7964w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7700w7963w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7779w7962w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7706w7971w7972w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7706w7971w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7544w7970w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7711w7979w7980w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7711w7979w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7548w7978w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7522w7987w7988w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7522w7987w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7550w7986w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7528w7995w7996w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7528w7995w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7552w7994w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7530w8003w8004w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7530w8003w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7554w8002w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7532w8011w8012w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7532w8011w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7556w8010w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7534w8019w8020w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7534w8019w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7558w8018w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7580w7803w7804w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7580w7803w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7719w7802w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7536w8027w8028w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7536w8027w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7560w8026w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7538w8035w8036w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7538w8035w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7562w8034w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7540w8043w8044w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7540w8043w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7564w8042w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7542w8051w8052w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7542w8051w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7566w8050w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7586w7811w7812w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7586w7811w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7722w7810w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7592w7819w7820w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7592w7819w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7725w7818w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7598w7827w7828w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7598w7827w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7728w7826w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7604w7835w7836w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7604w7835w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7731w7834w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7610w7843w7844w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7610w7843w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7734w7842w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7616w7851w7852w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7616w7851w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7737w7850w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7622w7859w7860w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7622w7859w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7740w7858w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8385w8592w8593w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8385w8592w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8524w8590w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8444w8674w8675w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8444w8674w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8553w8673w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8450w8682w8683w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8450w8682w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8556w8681w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8456w8690w8691w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8456w8690w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8559w8689w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8462w8698w8699w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8462w8698w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8562w8697w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8468w8706w8707w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8468w8706w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8565w8705w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8474w8714w8715w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8474w8714w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8568w8713w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8480w8722w8723w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8480w8722w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8571w8721w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8486w8730w8731w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8486w8730w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8574w8729w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8492w8738w8739w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8492w8738w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8577w8737w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8498w8746w8747w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8498w8746w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8580w8745w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8390w8602w8603w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8390w8602w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8526w8601w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8504w8754w8755w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8504w8754w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8583w8753w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8510w8762w8763w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8510w8762w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8586w8761w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8516w8770w8771w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8516w8770w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8358w8769w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8521w8778w8779w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8521w8778w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8362w8777w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8334w8786w8787w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8334w8786w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8364w8785w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8340w8794w8795w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8340w8794w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8366w8793w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8342w8802w8803w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8342w8802w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8368w8801w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8344w8810w8811w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8344w8810w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8370w8809w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8346w8818w8819w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8346w8818w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8372w8817w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8348w8826w8827w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8348w8826w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8374w8825w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8396w8610w8611w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8396w8610w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8529w8609w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8350w8834w8835w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8350w8834w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8376w8833w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8352w8842w8843w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8352w8842w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8378w8841w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8354w8850w8851w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8354w8850w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8380w8849w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8356w8858w8859w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8356w8858w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8382w8857w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8402w8618w8619w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8402w8618w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8532w8617w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8408w8626w8627w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8408w8626w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8535w8625w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8414w8634w8635w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8414w8634w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8538w8633w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8420w8642w8643w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8420w8642w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8541w8641w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8426w8650w8651w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8426w8650w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8544w8649w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8432w8658w8659w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8432w8658w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8547w8657w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8438w8666w8667w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8438w8666w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8550w8665w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9196w9394w9395w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9196w9394w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9329w9392w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9255w9476w9477w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9255w9476w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9358w9475w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9261w9484w9485w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9261w9484w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9361w9483w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9267w9492w9493w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9267w9492w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9364w9491w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9273w9500w9501w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9273w9500w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9367w9499w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9279w9508w9509w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9279w9508w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9370w9507w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9285w9516w9517w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9285w9516w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9373w9515w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9291w9524w9525w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9291w9524w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9376w9523w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9297w9532w9533w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9297w9532w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9379w9531w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9303w9540w9541w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9303w9540w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9382w9539w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9309w9548w9549w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9309w9548w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9385w9547w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9201w9404w9405w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9201w9404w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9331w9403w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9315w9556w9557w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9315w9556w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9388w9555w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9321w9564w9565w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9321w9564w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9167w9563w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9326w9572w9573w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9326w9572w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9171w9571w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9141w9580w9581w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9141w9580w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9173w9579w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9147w9588w9589w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9147w9588w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9175w9587w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9149w9596w9597w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9149w9596w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9177w9595w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9151w9604w9605w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9151w9604w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9179w9603w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9153w9612w9613w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9153w9612w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9181w9611w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9155w9620w9621w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9155w9620w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9183w9619w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9157w9628w9629w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9157w9628w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9185w9627w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9207w9412w9413w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9207w9412w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9334w9411w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9159w9636w9637w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9159w9636w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9187w9635w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9161w9644w9645w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9161w9644w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9189w9643w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9163w9652w9653w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9163w9652w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9191w9651w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9165w9660w9661w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9165w9660w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9193w9659w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9213w9420w9421w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9213w9420w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9337w9419w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9219w9428w9429w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9219w9428w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9340w9427w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9225w9436w9437w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9225w9436w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9343w9435w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9231w9444w9445w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9231w9444w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9346w9443w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9237w9452w9453w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9237w9452w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9349w9451w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9243w9460w9461w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9243w9460w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9352w9459w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9249w9468w9469w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9249w9468w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9355w9467w(0);
	wire_ccc_cordic_m_w10192w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10002w10191w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10129w10189w(0);
	wire_ccc_cordic_m_w10274w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10061w10273w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10158w10272w(0);
	wire_ccc_cordic_m_w10282w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10067w10281w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10161w10280w(0);
	wire_ccc_cordic_m_w10290w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10073w10289w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10164w10288w(0);
	wire_ccc_cordic_m_w10298w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10079w10297w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10167w10296w(0);
	wire_ccc_cordic_m_w10306w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10085w10305w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10170w10304w(0);
	wire_ccc_cordic_m_w10314w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10091w10313w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10173w10312w(0);
	wire_ccc_cordic_m_w10322w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10097w10321w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10176w10320w(0);
	wire_ccc_cordic_m_w10330w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10103w10329w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10179w10328w(0);
	wire_ccc_cordic_m_w10338w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10109w10337w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10182w10336w(0);
	wire_ccc_cordic_m_w10346w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10115w10345w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10185w10344w(0);
	wire_ccc_cordic_m_w10202w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10007w10201w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10131w10200w(0);
	wire_ccc_cordic_m_w10354w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10121w10353w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9971w10352w(0);
	wire_ccc_cordic_m_w10362w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10126w10361w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9975w10360w(0);
	wire_ccc_cordic_m_w10370w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9943w10369w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9977w10368w(0);
	wire_ccc_cordic_m_w10378w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9949w10377w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9979w10376w(0);
	wire_ccc_cordic_m_w10386w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9951w10385w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9981w10384w(0);
	wire_ccc_cordic_m_w10394w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9953w10393w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9983w10392w(0);
	wire_ccc_cordic_m_w10402w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9955w10401w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9985w10400w(0);
	wire_ccc_cordic_m_w10410w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9957w10409w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9987w10408w(0);
	wire_ccc_cordic_m_w10418w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9959w10417w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9989w10416w(0);
	wire_ccc_cordic_m_w10426w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9961w10425w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9991w10424w(0);
	wire_ccc_cordic_m_w10210w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10013w10209w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10134w10208w(0);
	wire_ccc_cordic_m_w10434w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9963w10433w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9993w10432w(0);
	wire_ccc_cordic_m_w10442w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9965w10441w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9995w10440w(0);
	wire_ccc_cordic_m_w10450w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9967w10449w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9997w10448w(0);
	wire_ccc_cordic_m_w10458w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9969w10457w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9999w10456w(0);
	wire_ccc_cordic_m_w10218w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10019w10217w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10137w10216w(0);
	wire_ccc_cordic_m_w10226w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10025w10225w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10140w10224w(0);
	wire_ccc_cordic_m_w10234w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10031w10233w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10143w10232w(0);
	wire_ccc_cordic_m_w10242w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10037w10241w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10146w10240w(0);
	wire_ccc_cordic_m_w10250w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10043w10249w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10149w10248w(0);
	wire_ccc_cordic_m_w10258w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10049w10257w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10152w10256w(0);
	wire_ccc_cordic_m_w10266w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10055w10265w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10155w10264w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range861w1149w1150w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range861w1149w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1054w1147w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range920w1231w1232w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range920w1231w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1083w1230w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range926w1239w1240w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range926w1239w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1086w1238w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range932w1247w1248w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range932w1247w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1089w1246w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range938w1255w1256w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range938w1255w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1092w1254w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range944w1263w1264w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range944w1263w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1095w1262w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range950w1271w1272w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range950w1271w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1098w1270w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range956w1279w1280w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range956w1279w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1101w1278w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range962w1287w1288w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range962w1287w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1104w1286w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range968w1295w1296w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range968w1295w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1107w1294w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range974w1303w1304w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range974w1303w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1110w1302w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range866w1159w1160w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range866w1159w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1056w1158w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range980w1311w1312w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range980w1311w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1113w1310w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range986w1319w1320w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range986w1319w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1116w1318w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range992w1327w1328w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range992w1327w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1119w1326w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range998w1335w1336w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range998w1335w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1122w1334w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1004w1343w1344w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1004w1343w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1125w1342w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1010w1351w1352w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1010w1351w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1128w1350w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1016w1359w1360w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1016w1359w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1131w1358w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1022w1367w1368w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1022w1367w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1134w1366w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1028w1375w1376w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1028w1375w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1137w1374w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1034w1383w1384w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1034w1383w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1140w1382w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range872w1167w1168w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range872w1167w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1059w1166w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1040w1391w1392w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1040w1391w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1143w1390w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1046w1399w1400w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1046w1399w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range852w1398w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1051w1407w1408w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1051w1407w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range856w1406w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range846w1415w1416w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range846w1415w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range858w1414w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range878w1175w1176w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range878w1175w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1062w1174w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range884w1183w1184w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range884w1183w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1065w1182w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range890w1191w1192w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range890w1191w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1068w1190w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range896w1199w1200w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range896w1199w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1071w1198w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range902w1207w1208w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range902w1207w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1074w1206w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range908w1215w1216w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range908w1215w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1077w1214w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range914w1223w1224w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range914w1223w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1080w1222w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1717w1996w1997w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1717w1996w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1904w1994w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1776w2078w2079w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1776w2078w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1933w2077w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1782w2086w2087w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1782w2086w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1936w2085w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1788w2094w2095w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1788w2094w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1939w2093w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1794w2102w2103w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1794w2102w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1942w2101w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1800w2110w2111w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1800w2110w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1945w2109w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1806w2118w2119w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1806w2118w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1948w2117w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1812w2126w2127w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1812w2126w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1951w2125w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1818w2134w2135w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1818w2134w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1954w2133w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1824w2142w2143w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1824w2142w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1957w2141w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1830w2150w2151w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1830w2150w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1960w2149w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1722w2006w2007w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1722w2006w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1906w2005w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1836w2158w2159w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1836w2158w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1963w2157w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1842w2166w2167w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1842w2166w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1966w2165w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1848w2174w2175w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1848w2174w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1969w2173w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1854w2182w2183w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1854w2182w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1972w2181w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1860w2190w2191w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1860w2190w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1975w2189w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1866w2198w2199w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1866w2198w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1978w2197w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1872w2206w2207w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1872w2206w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1981w2205w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1878w2214w2215w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1878w2214w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1984w2213w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1884w2222w2223w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1884w2222w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1987w2221w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1890w2230w2231w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1890w2230w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1990w2229w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1728w2014w2015w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1728w2014w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1909w2013w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1896w2238w2239w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1896w2238w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1706w2237w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1901w2246w2247w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1901w2246w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1710w2245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1698w2254w2255w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1698w2254w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1712w2253w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1704w2262w2263w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1704w2262w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1714w2261w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1734w2022w2023w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1734w2022w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1912w2021w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1740w2030w2031w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1740w2030w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1915w2029w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1746w2038w2039w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1746w2038w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1918w2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1752w2046w2047w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1752w2046w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1921w2045w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1758w2054w2055w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1758w2054w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1924w2053w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1764w2062w2063w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1764w2062w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1927w2061w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1770w2070w2071w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1770w2070w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1930w2069w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2568w2838w2839w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2568w2838w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2749w2836w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2627w2920w2921w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2627w2920w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2778w2919w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2633w2928w2929w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2633w2928w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2781w2927w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2639w2936w2937w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2639w2936w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2784w2935w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2645w2944w2945w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2645w2944w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2787w2943w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2651w2952w2953w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2651w2952w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2790w2951w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2657w2960w2961w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2657w2960w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2793w2959w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2663w2968w2969w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2663w2968w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2796w2967w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2669w2976w2977w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2669w2976w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2799w2975w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2675w2984w2985w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2675w2984w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2802w2983w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2681w2992w2993w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2681w2992w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2805w2991w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2573w2848w2849w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2573w2848w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2751w2847w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2687w3000w3001w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2687w3000w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2808w2999w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2693w3008w3009w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2693w3008w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2811w3007w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2699w3016w3017w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2699w3016w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2814w3015w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2705w3024w3025w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2705w3024w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2817w3023w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2711w3032w3033w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2711w3032w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2820w3031w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2717w3040w3041w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2717w3040w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2823w3039w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2723w3048w3049w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2723w3048w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2826w3047w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2729w3056w3057w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2729w3056w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2829w3055w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2735w3064w3065w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2735w3064w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2832w3063w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2741w3072w3073w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2741w3072w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2555w3071w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2579w2856w2857w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2579w2856w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2754w2855w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2746w3080w3081w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2746w3080w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2559w3079w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2545w3088w3089w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2545w3088w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2561w3087w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2551w3096w3097w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2551w3096w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2563w3095w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2553w3104w3105w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2553w3104w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2565w3103w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2585w2864w2865w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2585w2864w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2757w2863w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2591w2872w2873w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2591w2872w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2760w2871w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2597w2880w2881w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2597w2880w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2763w2879w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2603w2888w2889w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2603w2888w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2766w2887w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2609w2896w2897w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2609w2896w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2769w2895w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2615w2904w2905w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2615w2904w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2772w2903w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2621w2912w2913w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2621w2912w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2775w2911w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3414w3675w3676w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3414w3675w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3589w3673w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3473w3757w3758w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3473w3757w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3618w3756w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3479w3765w3766w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3479w3765w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3621w3764w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3485w3773w3774w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3485w3773w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3624w3772w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3491w3781w3782w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3491w3781w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3627w3780w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3497w3789w3790w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3497w3789w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3630w3788w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3503w3797w3798w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3503w3797w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3633w3796w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3509w3805w3806w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3509w3805w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3636w3804w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3515w3813w3814w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3515w3813w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3639w3812w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3521w3821w3822w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3521w3821w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3642w3820w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3527w3829w3830w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3527w3829w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3645w3828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3419w3685w3686w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3419w3685w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3591w3684w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3533w3837w3838w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3533w3837w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3648w3836w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3539w3845w3846w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3539w3845w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3651w3844w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3545w3853w3854w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3545w3853w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3654w3852w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3551w3861w3862w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3551w3861w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3657w3860w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3557w3869w3870w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3557w3869w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3660w3868w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3563w3877w3878w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3563w3877w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3663w3876w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3569w3885w3886w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3569w3885w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3666w3884w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3575w3893w3894w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3575w3893w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3669w3892w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3581w3901w3902w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3581w3901w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3399w3900w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3586w3909w3910w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3586w3909w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3403w3908w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3425w3693w3694w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3425w3693w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3594w3692w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3387w3917w3918w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3387w3917w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3405w3916w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3393w3925w3926w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3393w3925w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3407w3924w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3395w3933w3934w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3395w3933w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3409w3932w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3397w3941w3942w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3397w3941w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3411w3940w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3431w3701w3702w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3431w3701w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3597w3700w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3437w3709w3710w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3437w3709w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3600w3708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3443w3717w3718w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3443w3717w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3603w3716w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3449w3725w3726w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3449w3725w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3606w3724w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3455w3733w3734w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3455w3733w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3609w3732w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3461w3741w3742w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3461w3741w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3612w3740w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3467w3749w3750w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3467w3749w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3615w3748w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4255w4507w4508w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4255w4507w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4424w4505w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4314w4589w4590w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4314w4589w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4453w4588w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4320w4597w4598w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4320w4597w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4456w4596w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4326w4605w4606w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4326w4605w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4459w4604w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4332w4613w4614w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4332w4613w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4462w4612w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4338w4621w4622w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4338w4621w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4465w4620w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4344w4629w4630w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4344w4629w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4468w4628w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4350w4637w4638w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4350w4637w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4471w4636w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4356w4645w4646w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4356w4645w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4474w4644w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4362w4653w4654w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4362w4653w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4477w4652w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4368w4661w4662w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4368w4661w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4480w4660w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4260w4517w4518w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4260w4517w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4426w4516w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4374w4669w4670w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4374w4669w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4483w4668w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4380w4677w4678w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4380w4677w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4486w4676w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4386w4685w4686w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4386w4685w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4489w4684w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4392w4693w4694w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4392w4693w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4492w4692w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4398w4701w4702w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4398w4701w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4495w4700w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4404w4709w4710w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4404w4709w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4498w4708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4410w4717w4718w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4410w4717w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4501w4716w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4416w4725w4726w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4416w4725w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4238w4724w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4421w4733w4734w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4421w4733w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4242w4732w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4224w4741w4742w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4224w4741w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4244w4740w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4266w4525w4526w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4266w4525w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4429w4524w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4230w4749w4750w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4230w4749w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4246w4748w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4232w4757w4758w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4232w4757w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4248w4756w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4234w4765w4766w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4234w4765w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4250w4764w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4236w4773w4774w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4236w4773w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4252w4772w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4272w4533w4534w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4272w4533w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4432w4532w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4278w4541w4542w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4278w4541w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4435w4540w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4284w4549w4550w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4284w4549w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4438w4548w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4290w4557w4558w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4290w4557w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4441w4556w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4296w4565w4566w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4296w4565w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4444w4564w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4302w4573w4574w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4302w4573w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4447w4572w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4308w4581w4582w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4308w4581w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4450w4580w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5091w5334w5335w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5091w5334w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5254w5332w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5150w5416w5417w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5150w5416w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5283w5415w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5156w5424w5425w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5156w5424w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5286w5423w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5162w5432w5433w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5162w5432w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5289w5431w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5168w5440w5441w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5168w5440w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5292w5439w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5174w5448w5449w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5174w5448w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5295w5447w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5180w5456w5457w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5180w5456w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5298w5455w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5186w5464w5465w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5186w5464w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5301w5463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5192w5472w5473w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5192w5472w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5304w5471w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5198w5480w5481w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5198w5480w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5307w5479w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5204w5488w5489w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5204w5488w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5310w5487w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5096w5344w5345w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5096w5344w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5256w5343w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5210w5496w5497w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5210w5496w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5313w5495w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5216w5504w5505w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5216w5504w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5316w5503w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5222w5512w5513w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5222w5512w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5319w5511w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5228w5520w5521w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5228w5520w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5322w5519w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5234w5528w5529w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5234w5528w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5325w5527w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5240w5536w5537w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5240w5536w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5328w5535w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5246w5544w5545w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5246w5544w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5072w5543w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5251w5552w5553w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5251w5552w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5076w5551w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5056w5560w5561w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5056w5560w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5078w5559w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5062w5568w5569w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5062w5568w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5080w5567w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5102w5352w5353w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5102w5352w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5259w5351w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5064w5576w5577w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5064w5576w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5082w5575w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5066w5584w5585w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5066w5584w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5084w5583w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5068w5592w5593w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5068w5592w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5086w5591w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5070w5600w5601w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5070w5600w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5088w5599w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5108w5360w5361w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5108w5360w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5262w5359w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5114w5368w5369w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5114w5368w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5265w5367w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5120w5376w5377w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5120w5376w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5268w5375w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5126w5384w5385w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5126w5384w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5271w5383w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5132w5392w5393w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5132w5392w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5274w5391w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5138w5400w5401w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5138w5400w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5277w5399w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5144w5408w5409w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5144w5408w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5280w5407w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5922w6156w6157w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5922w6156w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6079w6154w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5981w6238w6239w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5981w6238w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6108w6237w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5987w6246w6247w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5987w6246w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6111w6245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5993w6254w6255w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5993w6254w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6114w6253w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5999w6262w6263w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5999w6262w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6117w6261w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6005w6270w6271w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6005w6270w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6120w6269w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6011w6278w6279w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6011w6278w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6123w6277w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6017w6286w6287w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6017w6286w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6126w6285w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6023w6294w6295w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6023w6294w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6129w6293w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6029w6302w6303w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6029w6302w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6132w6301w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6035w6310w6311w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6035w6310w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6135w6309w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5927w6166w6167w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5927w6166w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6081w6165w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6041w6318w6319w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6041w6318w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6138w6317w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6047w6326w6327w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6047w6326w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6141w6325w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6053w6334w6335w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6053w6334w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6144w6333w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6059w6342w6343w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6059w6342w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6147w6341w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6065w6350w6351w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6065w6350w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6150w6349w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6071w6358w6359w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6071w6358w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5901w6357w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6076w6366w6367w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6076w6366w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5905w6365w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5883w6374w6375w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5883w6374w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5907w6373w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5889w6382w6383w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5889w6382w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5909w6381w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5891w6390w6391w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5891w6390w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5911w6389w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5933w6174w6175w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5933w6174w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6084w6173w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5893w6398w6399w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5893w6398w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5913w6397w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5895w6406w6407w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5895w6406w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5915w6405w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5897w6414w6415w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5897w6414w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5917w6413w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5899w6422w6423w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5899w6422w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5919w6421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5939w6182w6183w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5939w6182w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6087w6181w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5945w6190w6191w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5945w6190w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6090w6189w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5951w6198w6199w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5951w6198w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6093w6197w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5957w6206w6207w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5957w6206w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6096w6205w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5963w6214w6215w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5963w6214w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6099w6213w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5969w6222w6223w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5969w6222w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6102w6221w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5975w6230w6231w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5975w6230w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6105w6229w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6748w6973w6974w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6748w6973w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6899w6971w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6807w7055w7056w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6807w7055w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6928w7054w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6813w7063w7064w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6813w7063w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6931w7062w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6819w7071w7072w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6819w7071w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6934w7070w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6825w7079w7080w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6825w7079w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6937w7078w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6831w7087w7088w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6831w7087w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6940w7086w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6837w7095w7096w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6837w7095w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6943w7094w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6843w7103w7104w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6843w7103w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6946w7102w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6849w7111w7112w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6849w7111w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6949w7110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6855w7119w7120w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6855w7119w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6952w7118w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6861w7127w7128w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6861w7127w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6955w7126w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6753w6983w6984w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6753w6983w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6901w6982w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6867w7135w7136w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6867w7135w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6958w7134w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6873w7143w7144w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6873w7143w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6961w7142w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6879w7151w7152w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6879w7151w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6964w7150w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6885w7159w7160w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6885w7159w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6967w7158w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6891w7167w7168w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6891w7167w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6725w7166w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6896w7175w7176w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6896w7175w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6729w7174w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6705w7183w7184w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6705w7183w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6731w7182w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6711w7191w7192w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6711w7191w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6733w7190w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6713w7199w7200w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6713w7199w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6735w7198w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6715w7207w7208w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6715w7207w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6737w7206w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6759w6991w6992w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6759w6991w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6904w6990w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6717w7215w7216w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6717w7215w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6739w7214w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6719w7223w7224w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6719w7223w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6741w7222w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6721w7231w7232w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6721w7231w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6743w7230w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6723w7239w7240w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6723w7239w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6745w7238w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6765w6999w7000w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6765w6999w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6907w6998w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6771w7007w7008w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6771w7007w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6910w7006w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6777w7015w7016w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6777w7015w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6913w7014w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6783w7023w7024w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6783w7023w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6916w7022w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6789w7031w7032w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6789w7031w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6919w7030w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6795w7039w7040w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6795w7039w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6922w7038w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6801w7047w7048w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6801w7047w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6925w7046w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7572w7790w7791w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7572w7790w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7715w7789w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7631w7871w7872w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7631w7871w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7744w7870w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7637w7879w7880w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7637w7879w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7747w7878w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7643w7887w7888w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7643w7887w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7750w7886w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7649w7895w7896w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7649w7895w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7753w7894w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7655w7903w7904w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7655w7903w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7756w7902w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7661w7911w7912w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7661w7911w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7759w7910w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7667w7919w7920w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7667w7919w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7762w7918w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7673w7927w7928w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7673w7927w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7765w7926w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7679w7935w7936w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7679w7935w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7768w7934w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7685w7943w7944w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7685w7943w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7771w7942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7577w7799w7800w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7577w7799w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7717w7798w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7691w7951w7952w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7691w7951w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7774w7950w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7697w7959w7960w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7697w7959w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7777w7958w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7703w7967w7968w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7703w7967w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7780w7966w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7709w7975w7976w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7709w7975w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7546w7974w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7712w7983w7984w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7712w7983w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7549w7982w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7526w7991w7992w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7526w7991w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7551w7990w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7529w7999w8000w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7529w7999w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7553w7998w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7531w8007w8008w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7531w8007w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7555w8006w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7533w8015w8016w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7533w8015w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7557w8014w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7535w8023w8024w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7535w8023w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7559w8022w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7583w7807w7808w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7583w7807w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7720w7806w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7537w8031w8032w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7537w8031w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7561w8030w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7539w8039w8040w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7539w8039w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7563w8038w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7541w8047w8048w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7541w8047w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7565w8046w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7543w8055w8056w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7543w8055w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7567w8054w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7589w7815w7816w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7589w7815w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7723w7814w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7595w7823w7824w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7595w7823w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7726w7822w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7601w7831w7832w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7601w7831w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7729w7830w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7607w7839w7840w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7607w7839w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7732w7838w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7613w7847w7848w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7613w7847w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7735w7846w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7619w7855w7856w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7619w7855w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7738w7854w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7625w7863w7864w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7625w7863w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7741w7862w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8388w8597w8598w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8388w8597w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8525w8596w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8447w8678w8679w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8447w8678w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8554w8677w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8453w8686w8687w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8453w8686w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8557w8685w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8459w8694w8695w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8459w8694w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8560w8693w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8465w8702w8703w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8465w8702w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8563w8701w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8471w8710w8711w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8471w8710w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8566w8709w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8477w8718w8719w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8477w8718w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8569w8717w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8483w8726w8727w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8483w8726w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8572w8725w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8489w8734w8735w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8489w8734w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8575w8733w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8495w8742w8743w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8495w8742w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8578w8741w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8501w8750w8751w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8501w8750w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8581w8749w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8393w8606w8607w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8393w8606w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8527w8605w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8507w8758w8759w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8507w8758w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8584w8757w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8513w8766w8767w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8513w8766w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8587w8765w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8519w8774w8775w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8519w8774w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8360w8773w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8522w8782w8783w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8522w8782w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8363w8781w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8338w8790w8791w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8338w8790w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8365w8789w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8341w8798w8799w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8341w8798w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8367w8797w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8343w8806w8807w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8343w8806w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8369w8805w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8345w8814w8815w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8345w8814w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8371w8813w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8347w8822w8823w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8347w8822w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8373w8821w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8349w8830w8831w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8349w8830w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8375w8829w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8399w8614w8615w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8399w8614w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8530w8613w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8351w8838w8839w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8351w8838w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8377w8837w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8353w8846w8847w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8353w8846w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8379w8845w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8355w8854w8855w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8355w8854w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8381w8853w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8357w8862w8863w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8357w8862w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8383w8861w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8405w8622w8623w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8405w8622w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8533w8621w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8411w8630w8631w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8411w8630w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8536w8629w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8417w8638w8639w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8417w8638w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8539w8637w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8423w8646w8647w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8423w8646w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8542w8645w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8429w8654w8655w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8429w8654w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8545w8653w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8435w8662w8663w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8435w8662w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8548w8661w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8441w8670w8671w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8441w8670w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8551w8669w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9199w9399w9400w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9199w9399w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9330w9398w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9258w9480w9481w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9258w9480w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9359w9479w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9264w9488w9489w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9264w9488w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9362w9487w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9270w9496w9497w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9270w9496w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9365w9495w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9276w9504w9505w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9276w9504w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9368w9503w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9282w9512w9513w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9282w9512w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9371w9511w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9288w9520w9521w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9288w9520w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9374w9519w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9294w9528w9529w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9294w9528w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9377w9527w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9300w9536w9537w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9300w9536w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9380w9535w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9306w9544w9545w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9306w9544w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9383w9543w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9312w9552w9553w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9312w9552w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9386w9551w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9204w9408w9409w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9204w9408w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9332w9407w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9318w9560w9561w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9318w9560w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9389w9559w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9324w9568w9569w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9324w9568w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9169w9567w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9327w9576w9577w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9327w9576w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9172w9575w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9145w9584w9585w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9145w9584w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9174w9583w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9148w9592w9593w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9148w9592w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9176w9591w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9150w9600w9601w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9150w9600w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9178w9599w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9152w9608w9609w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9152w9608w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9180w9607w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9154w9616w9617w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9154w9616w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9182w9615w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9156w9624w9625w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9156w9624w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9184w9623w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9158w9632w9633w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9158w9632w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9186w9631w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9210w9416w9417w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9210w9416w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9335w9415w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9160w9640w9641w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9160w9640w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9188w9639w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9162w9648w9649w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9162w9648w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9190w9647w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9164w9656w9657w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9164w9656w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9192w9655w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9166w9664w9665w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9166w9664w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9194w9663w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9216w9424w9425w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9216w9424w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9338w9423w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9222w9432w9433w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9222w9432w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9341w9431w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9228w9440w9441w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9228w9440w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9344w9439w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9234w9448w9449w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9234w9448w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9347w9447w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9240w9456w9457w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9240w9456w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9350w9455w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9246w9464w9465w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9246w9464w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9353w9463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9252w9472w9473w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9252w9472w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9356w9471w(0);
	wire_ccc_cordic_m_w10197w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10005w10196w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10130w10195w(0);
	wire_ccc_cordic_m_w10278w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10064w10277w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10159w10276w(0);
	wire_ccc_cordic_m_w10286w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10070w10285w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10162w10284w(0);
	wire_ccc_cordic_m_w10294w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10076w10293w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10165w10292w(0);
	wire_ccc_cordic_m_w10302w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10082w10301w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10168w10300w(0);
	wire_ccc_cordic_m_w10310w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10088w10309w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10171w10308w(0);
	wire_ccc_cordic_m_w10318w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10094w10317w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10174w10316w(0);
	wire_ccc_cordic_m_w10326w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10100w10325w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10177w10324w(0);
	wire_ccc_cordic_m_w10334w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10106w10333w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10180w10332w(0);
	wire_ccc_cordic_m_w10342w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10112w10341w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10183w10340w(0);
	wire_ccc_cordic_m_w10350w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10118w10349w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10186w10348w(0);
	wire_ccc_cordic_m_w10206w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10010w10205w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10132w10204w(0);
	wire_ccc_cordic_m_w10358w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10124w10357w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9973w10356w(0);
	wire_ccc_cordic_m_w10366w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10127w10365w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9976w10364w(0);
	wire_ccc_cordic_m_w10374w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9947w10373w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9978w10372w(0);
	wire_ccc_cordic_m_w10382w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9950w10381w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9980w10380w(0);
	wire_ccc_cordic_m_w10390w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9952w10389w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9982w10388w(0);
	wire_ccc_cordic_m_w10398w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9954w10397w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9984w10396w(0);
	wire_ccc_cordic_m_w10406w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9956w10405w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9986w10404w(0);
	wire_ccc_cordic_m_w10414w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9958w10413w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9988w10412w(0);
	wire_ccc_cordic_m_w10422w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9960w10421w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9990w10420w(0);
	wire_ccc_cordic_m_w10430w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9962w10429w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9992w10428w(0);
	wire_ccc_cordic_m_w10214w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10016w10213w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10135w10212w(0);
	wire_ccc_cordic_m_w10438w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9964w10437w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9994w10436w(0);
	wire_ccc_cordic_m_w10446w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9966w10445w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9996w10444w(0);
	wire_ccc_cordic_m_w10454w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9968w10453w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9998w10452w(0);
	wire_ccc_cordic_m_w10462w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9970w10461w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10000w10460w(0);
	wire_ccc_cordic_m_w10222w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10022w10221w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10138w10220w(0);
	wire_ccc_cordic_m_w10230w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10028w10229w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10141w10228w(0);
	wire_ccc_cordic_m_w10238w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10034w10237w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10144w10236w(0);
	wire_ccc_cordic_m_w10246w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10040w10245w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10147w10244w(0);
	wire_ccc_cordic_m_w10254w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10046w10253w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10150w10252w(0);
	wire_ccc_cordic_m_w10262w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10052w10261w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10153w10260w(0);
	wire_ccc_cordic_m_w10270w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10058w10269w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10156w10268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range864w1154w1155w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range864w1154w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1055w1153w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range923w1235w1236w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range923w1235w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1084w1234w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range929w1243w1244w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range929w1243w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1087w1242w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range935w1251w1252w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range935w1251w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1090w1250w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range941w1259w1260w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range941w1259w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1093w1258w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range947w1267w1268w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range947w1267w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1096w1266w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range953w1275w1276w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range953w1275w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1099w1274w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range959w1283w1284w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range959w1283w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1102w1282w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range965w1291w1292w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range965w1291w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1105w1290w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range971w1299w1300w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range971w1299w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1108w1298w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range977w1307w1308w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range977w1307w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1111w1306w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range869w1163w1164w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range869w1163w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1057w1162w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range983w1315w1316w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range983w1315w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1114w1314w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range989w1323w1324w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range989w1323w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1117w1322w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range995w1331w1332w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range995w1331w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1120w1330w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1001w1339w1340w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1001w1339w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1123w1338w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1007w1347w1348w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1007w1347w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1126w1346w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1013w1355w1356w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1013w1355w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1129w1354w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1019w1363w1364w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1019w1363w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1132w1362w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1025w1371w1372w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1025w1371w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1135w1370w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1031w1379w1380w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1031w1379w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1138w1378w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1037w1387w1388w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1037w1387w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1141w1386w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range875w1171w1172w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range875w1171w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1060w1170w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1043w1395w1396w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1043w1395w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1144w1394w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1049w1403w1404w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1049w1403w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range854w1402w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1052w1411w1412w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1052w1411w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range857w1410w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range850w1419w1420w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range850w1419w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range859w1418w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range881w1179w1180w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range881w1179w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1063w1178w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range887w1187w1188w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range887w1187w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1066w1186w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range893w1195w1196w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range893w1195w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1069w1194w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range899w1203w1204w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range899w1203w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1072w1202w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range905w1211w1212w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range905w1211w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1075w1210w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range911w1219w1220w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range911w1219w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1078w1218w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range917w1227w1228w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range917w1227w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1081w1226w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1720w2001w2002w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1720w2001w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1905w2000w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1779w2082w2083w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1779w2082w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1934w2081w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1785w2090w2091w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1785w2090w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1937w2089w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1791w2098w2099w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1791w2098w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1940w2097w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1797w2106w2107w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1797w2106w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1943w2105w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1803w2114w2115w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1803w2114w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1946w2113w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1809w2122w2123w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1809w2122w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1949w2121w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1815w2130w2131w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1815w2130w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1952w2129w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1821w2138w2139w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1821w2138w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1955w2137w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1827w2146w2147w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1827w2146w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1958w2145w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1833w2154w2155w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1833w2154w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1961w2153w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1725w2010w2011w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1725w2010w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1907w2009w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1839w2162w2163w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1839w2162w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1964w2161w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1845w2170w2171w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1845w2170w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1967w2169w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1851w2178w2179w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1851w2178w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1970w2177w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1857w2186w2187w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1857w2186w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1973w2185w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1863w2194w2195w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1863w2194w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1976w2193w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1869w2202w2203w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1869w2202w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1979w2201w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1875w2210w2211w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1875w2210w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1982w2209w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1881w2218w2219w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1881w2218w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1985w2217w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1887w2226w2227w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1887w2226w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1988w2225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1893w2234w2235w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1893w2234w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1991w2233w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1731w2018w2019w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1731w2018w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1910w2017w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1899w2242w2243w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1899w2242w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1708w2241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1902w2250w2251w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1902w2250w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1711w2249w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1702w2258w2259w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1702w2258w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1713w2257w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1705w2266w2267w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1705w2266w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1715w2265w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1737w2026w2027w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1737w2026w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1913w2025w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1743w2034w2035w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1743w2034w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1916w2033w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1749w2042w2043w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1749w2042w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1919w2041w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1755w2050w2051w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1755w2050w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1922w2049w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1761w2058w2059w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1761w2058w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1925w2057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1767w2066w2067w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1767w2066w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1928w2065w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1773w2074w2075w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1773w2074w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1931w2073w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2571w2843w2844w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2571w2843w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2750w2842w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2630w2924w2925w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2630w2924w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2779w2923w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2636w2932w2933w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2636w2932w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2782w2931w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2642w2940w2941w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2642w2940w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2785w2939w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2648w2948w2949w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2648w2948w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2788w2947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2654w2956w2957w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2654w2956w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2791w2955w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2660w2964w2965w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2660w2964w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2794w2963w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2666w2972w2973w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2666w2972w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2797w2971w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2672w2980w2981w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2672w2980w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2800w2979w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2678w2988w2989w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2678w2988w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2803w2987w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2684w2996w2997w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2684w2996w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2806w2995w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2576w2852w2853w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2576w2852w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2752w2851w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2690w3004w3005w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2690w3004w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2809w3003w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2696w3012w3013w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2696w3012w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2812w3011w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2702w3020w3021w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2702w3020w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2815w3019w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2708w3028w3029w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2708w3028w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2818w3027w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2714w3036w3037w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2714w3036w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2821w3035w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2720w3044w3045w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2720w3044w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2824w3043w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2726w3052w3053w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2726w3052w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2827w3051w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2732w3060w3061w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2732w3060w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2830w3059w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2738w3068w3069w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2738w3068w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2833w3067w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2744w3076w3077w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2744w3076w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2557w3075w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2582w2860w2861w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2582w2860w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2755w2859w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2747w3084w3085w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2747w3084w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2560w3083w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2549w3092w3093w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2549w3092w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2562w3091w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2552w3100w3101w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2552w3100w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2564w3099w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2554w3108w3109w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2554w3108w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2566w3107w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2588w2868w2869w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2588w2868w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2758w2867w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2594w2876w2877w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2594w2876w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2761w2875w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2600w2884w2885w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2600w2884w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2764w2883w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2606w2892w2893w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2606w2892w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2767w2891w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2612w2900w2901w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2612w2900w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2770w2899w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2618w2908w2909w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2618w2908w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2773w2907w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2624w2916w2917w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2624w2916w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2776w2915w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3417w3680w3681w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3417w3680w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3590w3679w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3476w3761w3762w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3476w3761w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3619w3760w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3482w3769w3770w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3482w3769w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3622w3768w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3488w3777w3778w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3488w3777w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3625w3776w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3494w3785w3786w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3494w3785w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3628w3784w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3500w3793w3794w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3500w3793w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3631w3792w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3506w3801w3802w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3506w3801w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3634w3800w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3512w3809w3810w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3512w3809w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3637w3808w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3518w3817w3818w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3518w3817w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3640w3816w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3524w3825w3826w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3524w3825w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3643w3824w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3530w3833w3834w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3530w3833w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3646w3832w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3422w3689w3690w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3422w3689w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3592w3688w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3536w3841w3842w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3536w3841w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3649w3840w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3542w3849w3850w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3542w3849w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3652w3848w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3548w3857w3858w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3548w3857w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3655w3856w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3554w3865w3866w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3554w3865w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3658w3864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3560w3873w3874w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3560w3873w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3661w3872w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3566w3881w3882w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3566w3881w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3664w3880w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3572w3889w3890w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3572w3889w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3667w3888w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3578w3897w3898w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3578w3897w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3670w3896w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3584w3905w3906w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3584w3905w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3401w3904w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3587w3913w3914w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3587w3913w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3404w3912w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3428w3697w3698w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3428w3697w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3595w3696w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3391w3921w3922w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3391w3921w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3406w3920w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3394w3929w3930w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3394w3929w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3408w3928w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3396w3937w3938w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3396w3937w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3410w3936w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3398w3945w3946w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3398w3945w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3412w3944w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3434w3705w3706w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3434w3705w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3598w3704w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3440w3713w3714w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3440w3713w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3601w3712w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3446w3721w3722w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3446w3721w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3604w3720w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3452w3729w3730w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3452w3729w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3607w3728w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3458w3737w3738w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3458w3737w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3610w3736w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3464w3745w3746w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3464w3745w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3613w3744w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3470w3753w3754w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3470w3753w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3616w3752w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4258w4512w4513w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4258w4512w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4425w4511w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4317w4593w4594w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4317w4593w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4454w4592w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4323w4601w4602w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4323w4601w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4457w4600w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4329w4609w4610w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4329w4609w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4460w4608w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4335w4617w4618w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4335w4617w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4463w4616w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4341w4625w4626w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4341w4625w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4466w4624w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4347w4633w4634w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4347w4633w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4469w4632w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4353w4641w4642w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4353w4641w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4472w4640w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4359w4649w4650w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4359w4649w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4475w4648w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4365w4657w4658w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4365w4657w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4478w4656w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4371w4665w4666w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4371w4665w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4481w4664w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4263w4521w4522w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4263w4521w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4427w4520w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4377w4673w4674w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4377w4673w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4484w4672w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4383w4681w4682w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4383w4681w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4487w4680w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4389w4689w4690w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4389w4689w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4490w4688w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4395w4697w4698w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4395w4697w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4493w4696w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4401w4705w4706w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4401w4705w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4496w4704w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4407w4713w4714w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4407w4713w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4499w4712w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4413w4721w4722w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4413w4721w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4502w4720w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4419w4729w4730w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4419w4729w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4240w4728w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4422w4737w4738w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4422w4737w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4243w4736w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4228w4745w4746w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4228w4745w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4245w4744w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4269w4529w4530w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4269w4529w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4430w4528w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4231w4753w4754w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4231w4753w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4247w4752w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4233w4761w4762w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4233w4761w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4249w4760w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4235w4769w4770w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4235w4769w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4251w4768w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4237w4777w4778w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4237w4777w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4253w4776w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4275w4537w4538w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4275w4537w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4433w4536w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4281w4545w4546w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4281w4545w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4436w4544w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4287w4553w4554w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4287w4553w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4439w4552w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4293w4561w4562w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4293w4561w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4442w4560w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4299w4569w4570w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4299w4569w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4445w4568w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4305w4577w4578w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4305w4577w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4448w4576w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4311w4585w4586w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4311w4585w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4451w4584w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5094w5339w5340w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5094w5339w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5255w5338w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5153w5420w5421w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5153w5420w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5284w5419w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5159w5428w5429w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5159w5428w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5287w5427w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5165w5436w5437w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5165w5436w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5290w5435w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5171w5444w5445w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5171w5444w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5293w5443w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5177w5452w5453w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5177w5452w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5296w5451w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5183w5460w5461w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5183w5460w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5299w5459w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5189w5468w5469w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5189w5468w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5302w5467w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5195w5476w5477w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5195w5476w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5305w5475w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5201w5484w5485w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5201w5484w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5308w5483w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5207w5492w5493w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5207w5492w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5311w5491w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5099w5348w5349w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5099w5348w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5257w5347w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5213w5500w5501w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5213w5500w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5314w5499w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5219w5508w5509w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5219w5508w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5317w5507w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5225w5516w5517w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5225w5516w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5320w5515w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5231w5524w5525w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5231w5524w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5323w5523w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5237w5532w5533w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5237w5532w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5326w5531w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5243w5540w5541w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5243w5540w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5329w5539w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5249w5548w5549w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5249w5548w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5074w5547w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5252w5556w5557w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5252w5556w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5077w5555w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5060w5564w5565w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5060w5564w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5079w5563w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5063w5572w5573w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5063w5572w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5081w5571w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5105w5356w5357w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5105w5356w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5260w5355w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5065w5580w5581w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5065w5580w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5083w5579w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5067w5588w5589w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5067w5588w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5085w5587w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5069w5596w5597w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5069w5596w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5087w5595w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5071w5604w5605w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5071w5604w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5089w5603w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5111w5364w5365w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5111w5364w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5263w5363w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5117w5372w5373w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5117w5372w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5266w5371w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5123w5380w5381w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5123w5380w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5269w5379w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5129w5388w5389w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5129w5388w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5272w5387w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5135w5396w5397w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5135w5396w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5275w5395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5141w5404w5405w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5141w5404w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5278w5403w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5147w5412w5413w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5147w5412w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5281w5411w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5925w6161w6162w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5925w6161w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6080w6160w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5984w6242w6243w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5984w6242w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6109w6241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5990w6250w6251w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5990w6250w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6112w6249w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5996w6258w6259w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5996w6258w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6115w6257w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6002w6266w6267w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6002w6266w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6118w6265w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6008w6274w6275w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6008w6274w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6121w6273w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6014w6282w6283w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6014w6282w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6124w6281w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6020w6290w6291w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6020w6290w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6127w6289w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6026w6298w6299w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6026w6298w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6130w6297w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6032w6306w6307w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6032w6306w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6133w6305w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6038w6314w6315w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6038w6314w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6136w6313w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5930w6170w6171w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5930w6170w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6082w6169w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6044w6322w6323w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6044w6322w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6139w6321w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6050w6330w6331w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6050w6330w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6142w6329w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6056w6338w6339w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6056w6338w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6145w6337w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6062w6346w6347w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6062w6346w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6148w6345w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6068w6354w6355w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6068w6354w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6151w6353w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6074w6362w6363w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6074w6362w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5903w6361w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6077w6370w6371w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6077w6370w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5906w6369w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5887w6378w6379w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5887w6378w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5908w6377w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5890w6386w6387w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5890w6386w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5910w6385w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5892w6394w6395w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5892w6394w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5912w6393w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5936w6178w6179w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5936w6178w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6085w6177w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5894w6402w6403w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5894w6402w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5914w6401w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5896w6410w6411w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5896w6410w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5916w6409w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5898w6418w6419w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5898w6418w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5918w6417w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5900w6426w6427w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5900w6426w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5920w6425w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5942w6186w6187w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5942w6186w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6088w6185w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5948w6194w6195w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5948w6194w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6091w6193w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5954w6202w6203w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5954w6202w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6094w6201w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5960w6210w6211w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5960w6210w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6097w6209w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5966w6218w6219w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5966w6218w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6100w6217w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5972w6226w6227w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5972w6226w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6103w6225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5978w6234w6235w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5978w6234w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6106w6233w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6751w6978w6979w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6751w6978w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6900w6977w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6810w7059w7060w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6810w7059w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6929w7058w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6816w7067w7068w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6816w7067w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6932w7066w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6822w7075w7076w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6822w7075w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6935w7074w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6828w7083w7084w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6828w7083w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6938w7082w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6834w7091w7092w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6834w7091w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6941w7090w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6840w7099w7100w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6840w7099w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6944w7098w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6846w7107w7108w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6846w7107w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6947w7106w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6852w7115w7116w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6852w7115w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6950w7114w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6858w7123w7124w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6858w7123w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6953w7122w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6864w7131w7132w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6864w7131w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6956w7130w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6756w6987w6988w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6756w6987w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6902w6986w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6870w7139w7140w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6870w7139w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6959w7138w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6876w7147w7148w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6876w7147w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6962w7146w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6882w7155w7156w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6882w7155w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6965w7154w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6888w7163w7164w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6888w7163w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6968w7162w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6894w7171w7172w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6894w7171w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6727w7170w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6897w7179w7180w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6897w7179w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6730w7178w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6709w7187w7188w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6709w7187w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6732w7186w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6712w7195w7196w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6712w7195w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6734w7194w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6714w7203w7204w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6714w7203w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6736w7202w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6716w7211w7212w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6716w7211w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6738w7210w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6762w6995w6996w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6762w6995w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6905w6994w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6718w7219w7220w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6718w7219w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6740w7218w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6720w7227w7228w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6720w7227w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6742w7226w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6722w7235w7236w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6722w7235w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6744w7234w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6724w7243w7244w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6724w7243w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6746w7242w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6768w7003w7004w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6768w7003w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6908w7002w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6774w7011w7012w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6774w7011w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6911w7010w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6780w7019w7020w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6780w7019w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6914w7018w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6786w7027w7028w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6786w7027w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6917w7026w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6792w7035w7036w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6792w7035w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6920w7034w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6798w7043w7044w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6798w7043w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6923w7042w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6804w7051w7052w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6804w7051w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6926w7050w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8871w8873w8874w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8871w8873w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8952w8954w8955w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8952w8954w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8960w8962w8963w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8960w8962w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8968w8970w8971w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8968w8970w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8976w8978w8979w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8976w8978w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8984w8986w8987w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8984w8986w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8992w8994w8995w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8992w8994w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9000w9002w9003w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9000w9002w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9008w9010w9011w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9008w9010w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9016w9018w9019w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9016w9018w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9024w9026w9027w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9024w9026w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8880w8882w8883w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8880w8882w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9032w9034w9035w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9032w9034w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9040w9042w9043w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9040w9042w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9048w9050w9051w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9048w9050w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9056w9058w9059w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9056w9058w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9064w9066w9067w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9064w9066w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9072w9074w9075w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9072w9074w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9080w9082w9083w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9080w9082w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9088w9090w9091w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9088w9090w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9096w9098w9099w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9096w9098w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9104w9106w9107w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9104w9106w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8888w8890w8891w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8888w8890w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9112w9114w9115w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9112w9114w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9120w9122w9123w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9120w9122w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9128w9130w9131w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9128w9130w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9136w9138w9139w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9136w9138w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8896w8898w8899w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8896w8898w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8904w8906w8907w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8904w8906w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8912w8914w8915w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8912w8914w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8920w8922w8923w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8920w8922w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8928w8930w8931w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8928w8930w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8936w8938w8939w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8936w8938w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8944w8946w8947w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8944w8946w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9673w9675w9676w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9673w9675w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9754w9756w9757w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9754w9756w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9762w9764w9765w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9762w9764w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9770w9772w9773w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9770w9772w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9778w9780w9781w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9778w9780w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9786w9788w9789w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9786w9788w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9794w9796w9797w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9794w9796w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9802w9804w9805w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9802w9804w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9810w9812w9813w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9810w9812w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9818w9820w9821w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9818w9820w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9826w9828w9829w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9826w9828w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9682w9684w9685w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9682w9684w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9834w9836w9837w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9834w9836w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9842w9844w9845w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9842w9844w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9850w9852w9853w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9850w9852w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9858w9860w9861w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9858w9860w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9866w9868w9869w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9866w9868w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9874w9876w9877w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9874w9876w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9882w9884w9885w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9882w9884w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9890w9892w9893w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9890w9892w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9898w9900w9901w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9898w9900w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9906w9908w9909w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9906w9908w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9690w9692w9693w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9690w9692w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9914w9916w9917w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9914w9916w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9922w9924w9925w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9922w9924w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9930w9932w9933w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9930w9932w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9938w9940w9941w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9938w9940w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9698w9700w9701w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9698w9700w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9706w9708w9709w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9706w9708w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9714w9716w9717w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9714w9716w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9722w9724w9725w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9722w9724w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9730w9732w9733w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9730w9732w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9738w9740w9741w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9738w9740w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9746w9748w9749w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9746w9748w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10470w10472w10473w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10470w10472w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10551w10553w10554w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10551w10553w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10559w10561w10562w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10559w10561w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10567w10569w10570w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10567w10569w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10575w10577w10578w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10575w10577w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10583w10585w10586w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10583w10585w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10591w10593w10594w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10591w10593w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10599w10601w10602w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10599w10601w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10607w10609w10610w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10607w10609w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10615w10617w10618w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10615w10617w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10623w10625w10626w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10623w10625w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10479w10481w10482w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10479w10481w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10631w10633w10634w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10631w10633w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10639w10641w10642w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10639w10641w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10647w10649w10650w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10647w10649w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10655w10657w10658w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10655w10657w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10663w10665w10666w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10663w10665w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10671w10673w10674w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10671w10673w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10679w10681w10682w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10679w10681w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10687w10689w10690w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10687w10689w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10695w10697w10698w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10695w10697w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10703w10705w10706w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10703w10705w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10487w10489w10490w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10487w10489w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10711w10713w10714w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10711w10713w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10719w10721w10722w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10719w10721w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10727w10729w10730w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10727w10729w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10735w10737w10738w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10735w10737w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10495w10497w10498w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10495w10497w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10503w10505w10506w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10503w10505w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10511w10513w10514w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10511w10513w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10519w10521w10522w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10519w10521w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10527w10529w10530w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10527w10529w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10535w10537w10538w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10535w10537w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10543w10545w10546w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10543w10545w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1428w1430w1431w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1428w1430w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1509w1511w1512w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1509w1511w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1517w1519w1520w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1517w1519w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1525w1527w1528w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1525w1527w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1533w1535w1536w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1533w1535w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1541w1543w1544w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1541w1543w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1549w1551w1552w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1549w1551w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1557w1559w1560w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1557w1559w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1565w1567w1568w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1565w1567w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1573w1575w1576w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1573w1575w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1581w1583w1584w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1581w1583w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1437w1439w1440w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1437w1439w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1589w1591w1592w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1589w1591w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1597w1599w1600w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1597w1599w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1605w1607w1608w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1605w1607w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1613w1615w1616w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1613w1615w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1621w1623w1624w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1621w1623w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1629w1631w1632w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1629w1631w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1637w1639w1640w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1637w1639w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1645w1647w1648w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1645w1647w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1653w1655w1656w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1653w1655w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1661w1663w1664w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1661w1663w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1445w1447w1448w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1445w1447w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1669w1671w1672w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1669w1671w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1677w1679w1680w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1677w1679w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1685w1687w1688w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1685w1687w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1693w1695w1696w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1693w1695w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1453w1455w1456w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1453w1455w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1461w1463w1464w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1461w1463w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1469w1471w1472w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1469w1471w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1477w1479w1480w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1477w1479w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1485w1487w1488w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1485w1487w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1493w1495w1496w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1493w1495w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1501w1503w1504w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1501w1503w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2275w2277w2278w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2275w2277w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2356w2358w2359w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2356w2358w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2364w2366w2367w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2364w2366w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2372w2374w2375w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2372w2374w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2380w2382w2383w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2380w2382w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2388w2390w2391w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2388w2390w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2396w2398w2399w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2396w2398w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2404w2406w2407w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2404w2406w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2412w2414w2415w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2412w2414w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2420w2422w2423w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2420w2422w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2428w2430w2431w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2428w2430w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2284w2286w2287w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2284w2286w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2436w2438w2439w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2436w2438w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2444w2446w2447w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2444w2446w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2452w2454w2455w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2452w2454w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2460w2462w2463w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2460w2462w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2468w2470w2471w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2468w2470w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2476w2478w2479w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2476w2478w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2484w2486w2487w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2484w2486w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2492w2494w2495w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2492w2494w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2500w2502w2503w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2500w2502w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2508w2510w2511w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2508w2510w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2292w2294w2295w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2292w2294w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2516w2518w2519w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2516w2518w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2524w2526w2527w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2524w2526w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2532w2534w2535w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2532w2534w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2540w2542w2543w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2540w2542w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2300w2302w2303w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2300w2302w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2308w2310w2311w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2308w2310w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2316w2318w2319w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2316w2318w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2324w2326w2327w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2324w2326w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2332w2334w2335w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2332w2334w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2340w2342w2343w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2340w2342w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2348w2350w2351w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2348w2350w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3117w3119w3120w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3117w3119w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3198w3200w3201w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3198w3200w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3206w3208w3209w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3206w3208w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3214w3216w3217w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3214w3216w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3222w3224w3225w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3222w3224w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3230w3232w3233w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3230w3232w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3238w3240w3241w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3238w3240w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3246w3248w3249w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3246w3248w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3254w3256w3257w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3254w3256w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3262w3264w3265w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3262w3264w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3270w3272w3273w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3270w3272w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3126w3128w3129w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3126w3128w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3278w3280w3281w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3278w3280w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3286w3288w3289w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3286w3288w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3294w3296w3297w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3294w3296w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3302w3304w3305w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3302w3304w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3310w3312w3313w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3310w3312w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3318w3320w3321w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3318w3320w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3326w3328w3329w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3326w3328w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3334w3336w3337w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3334w3336w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3342w3344w3345w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3342w3344w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3350w3352w3353w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3350w3352w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3134w3136w3137w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3134w3136w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3358w3360w3361w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3358w3360w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3366w3368w3369w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3366w3368w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3374w3376w3377w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3374w3376w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3382w3384w3385w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3382w3384w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3142w3144w3145w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3142w3144w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3150w3152w3153w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3150w3152w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3158w3160w3161w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3158w3160w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3166w3168w3169w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3166w3168w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3174w3176w3177w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3174w3176w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3182w3184w3185w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3182w3184w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3190w3192w3193w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3190w3192w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3954w3956w3957w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3954w3956w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4035w4037w4038w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4035w4037w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4043w4045w4046w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4043w4045w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4051w4053w4054w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4051w4053w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4059w4061w4062w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4059w4061w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4067w4069w4070w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4067w4069w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4075w4077w4078w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4075w4077w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4083w4085w4086w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4083w4085w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4091w4093w4094w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4091w4093w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4099w4101w4102w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4099w4101w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4107w4109w4110w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4107w4109w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3963w3965w3966w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3963w3965w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4115w4117w4118w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4115w4117w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4123w4125w4126w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4123w4125w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4131w4133w4134w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4131w4133w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4139w4141w4142w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4139w4141w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4147w4149w4150w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4147w4149w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4155w4157w4158w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4155w4157w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4163w4165w4166w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4163w4165w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4171w4173w4174w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4171w4173w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4179w4181w4182w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4179w4181w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4187w4189w4190w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4187w4189w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3971w3973w3974w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3971w3973w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4195w4197w4198w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4195w4197w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4203w4205w4206w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4203w4205w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4211w4213w4214w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4211w4213w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4219w4221w4222w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4219w4221w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3979w3981w3982w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3979w3981w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3987w3989w3990w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3987w3989w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3995w3997w3998w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3995w3997w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4003w4005w4006w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4003w4005w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4011w4013w4014w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4011w4013w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4019w4021w4022w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4019w4021w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4027w4029w4030w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4027w4029w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4786w4788w4789w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4786w4788w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4867w4869w4870w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4867w4869w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4875w4877w4878w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4875w4877w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4883w4885w4886w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4883w4885w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4891w4893w4894w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4891w4893w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4899w4901w4902w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4899w4901w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4907w4909w4910w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4907w4909w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4915w4917w4918w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4915w4917w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4923w4925w4926w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4923w4925w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4931w4933w4934w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4931w4933w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4939w4941w4942w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4939w4941w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4795w4797w4798w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4795w4797w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4947w4949w4950w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4947w4949w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4955w4957w4958w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4955w4957w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4963w4965w4966w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4963w4965w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4971w4973w4974w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4971w4973w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4979w4981w4982w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4979w4981w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4987w4989w4990w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4987w4989w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4995w4997w4998w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4995w4997w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5003w5005w5006w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5003w5005w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5011w5013w5014w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5011w5013w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5019w5021w5022w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5019w5021w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4803w4805w4806w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4803w4805w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5027w5029w5030w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5027w5029w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5035w5037w5038w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5035w5037w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5043w5045w5046w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5043w5045w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5051w5053w5054w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5051w5053w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4811w4813w4814w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4811w4813w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4819w4821w4822w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4819w4821w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4827w4829w4830w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4827w4829w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4835w4837w4838w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4835w4837w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4843w4845w4846w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4843w4845w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4851w4853w4854w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4851w4853w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4859w4861w4862w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4859w4861w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5613w5615w5616w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5613w5615w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5694w5696w5697w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5694w5696w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5702w5704w5705w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5702w5704w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5710w5712w5713w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5710w5712w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5718w5720w5721w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5718w5720w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5726w5728w5729w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5726w5728w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5734w5736w5737w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5734w5736w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5742w5744w5745w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5742w5744w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5750w5752w5753w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5750w5752w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5758w5760w5761w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5758w5760w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5766w5768w5769w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5766w5768w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5622w5624w5625w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5622w5624w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5774w5776w5777w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5774w5776w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5782w5784w5785w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5782w5784w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5790w5792w5793w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5790w5792w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5798w5800w5801w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5798w5800w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5806w5808w5809w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5806w5808w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5814w5816w5817w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5814w5816w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5822w5824w5825w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5822w5824w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5830w5832w5833w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5830w5832w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5838w5840w5841w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5838w5840w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5846w5848w5849w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5846w5848w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5630w5632w5633w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5630w5632w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5854w5856w5857w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5854w5856w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5862w5864w5865w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5862w5864w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5870w5872w5873w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5870w5872w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5878w5880w5881w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5878w5880w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5638w5640w5641w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5638w5640w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5646w5648w5649w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5646w5648w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5654w5656w5657w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5654w5656w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5662w5664w5665w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5662w5664w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5670w5672w5673w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5670w5672w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5678w5680w5681w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5678w5680w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5686w5688w5689w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5686w5688w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6435w6437w6438w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6435w6437w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6516w6518w6519w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6516w6518w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6524w6526w6527w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6524w6526w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6532w6534w6535w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6532w6534w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6540w6542w6543w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6540w6542w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6548w6550w6551w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6548w6550w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6556w6558w6559w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6556w6558w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6564w6566w6567w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6564w6566w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6572w6574w6575w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6572w6574w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6580w6582w6583w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6580w6582w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6588w6590w6591w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6588w6590w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6444w6446w6447w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6444w6446w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6596w6598w6599w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6596w6598w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6604w6606w6607w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6604w6606w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6612w6614w6615w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6612w6614w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6620w6622w6623w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6620w6622w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6628w6630w6631w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6628w6630w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6636w6638w6639w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6636w6638w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6644w6646w6647w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6644w6646w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6652w6654w6655w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6652w6654w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6660w6662w6663w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6660w6662w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6668w6670w6671w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6668w6670w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6452w6454w6455w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6452w6454w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6676w6678w6679w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6676w6678w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6684w6686w6687w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6684w6686w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6692w6694w6695w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6692w6694w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6700w6702w6703w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6700w6702w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6460w6462w6463w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6460w6462w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6468w6470w6471w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6468w6470w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6476w6478w6479w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6476w6478w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6484w6486w6487w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6484w6486w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6492w6494w6495w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6492w6494w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6500w6502w6503w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6500w6502w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6508w6510w6511w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6508w6510w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7252w7254w7255w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7252w7254w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7333w7335w7336w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7333w7335w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7341w7343w7344w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7341w7343w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7349w7351w7352w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7349w7351w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7357w7359w7360w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7357w7359w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7365w7367w7368w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7365w7367w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7373w7375w7376w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7373w7375w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7381w7383w7384w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7381w7383w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7389w7391w7392w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7389w7391w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7397w7399w7400w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7397w7399w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7405w7407w7408w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7405w7407w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7261w7263w7264w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7261w7263w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7413w7415w7416w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7413w7415w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7421w7423w7424w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7421w7423w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7429w7431w7432w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7429w7431w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7437w7439w7440w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7437w7439w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7445w7447w7448w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7445w7447w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7453w7455w7456w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7453w7455w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7461w7463w7464w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7461w7463w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7469w7471w7472w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7469w7471w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7477w7479w7480w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7477w7479w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7485w7487w7488w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7485w7487w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7269w7271w7272w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7269w7271w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7493w7495w7496w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7493w7495w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7501w7503w7504w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7501w7503w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7509w7511w7512w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7509w7511w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7517w7519w7520w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7517w7519w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7277w7279w7280w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7277w7279w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7285w7287w7288w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7285w7287w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7293w7295w7296w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7293w7295w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7301w7303w7304w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7301w7303w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7309w7311w7312w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7309w7311w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7317w7319w7320w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7317w7319w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7325w7327w7328w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7325w7327w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8064w8066w8067w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8064w8066w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8145w8147w8148w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8145w8147w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8153w8155w8156w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8153w8155w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8161w8163w8164w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8161w8163w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8169w8171w8172w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8169w8171w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8177w8179w8180w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8177w8179w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8185w8187w8188w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8185w8187w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8193w8195w8196w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8193w8195w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8201w8203w8204w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8201w8203w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8209w8211w8212w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8209w8211w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8217w8219w8220w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8217w8219w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8073w8075w8076w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8073w8075w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8225w8227w8228w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8225w8227w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8233w8235w8236w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8233w8235w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8241w8243w8244w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8241w8243w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8249w8251w8252w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8249w8251w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8257w8259w8260w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8257w8259w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8265w8267w8268w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8265w8267w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8273w8275w8276w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8273w8275w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8281w8283w8284w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8281w8283w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8289w8291w8292w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8289w8291w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8297w8299w8300w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8297w8299w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8081w8083w8084w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8081w8083w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8305w8307w8308w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8305w8307w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8313w8315w8316w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8313w8315w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8321w8323w8324w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8321w8323w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8329w8331w8332w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8329w8331w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8089w8091w8092w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8089w8091w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8097w8099w8100w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8097w8099w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8105w8107w8108w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8105w8107w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8113w8115w8116w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8113w8115w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8121w8123w8124w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8121w8123w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8129w8131w8132w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8129w8131w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8137w8139w8140w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8137w8139w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	loop31 : FOR i IN 0 TO 33 GENERATE 
		wire_ccc_cordic_m_w_lg_estimate_w10920w(i) <= estimate_w(i) XOR wire_sincosbitff_w_lg_w_q_range10746w10747w(0);
	END GENERATE loop31;
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7782w8059w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7782w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7865w8142w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7865w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7873w8150w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7873w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7881w8158w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7881w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7889w8166w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7889w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7897w8174w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7897w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7905w8182w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7905w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7913w8190w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7913w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7921w8198w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7921w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7929w8206w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7929w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7937w8214w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7937w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7793w8070w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7793w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7945w8222w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7945w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7953w8230w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7953w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7961w8238w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7961w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7969w8246w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7969w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7977w8254w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7977w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7985w8262w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7985w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7993w8270w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7993w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8001w8278w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range8001w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8009w8286w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range8009w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8017w8294w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range8017w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7801w8078w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7801w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8025w8302w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range8025w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8033w8310w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range8033w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8041w8318w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range8041w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8049w8326w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range8049w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7809w8086w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7809w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7817w8094w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7817w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7825w8102w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7825w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7833w8110w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7833w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7841w8118w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7841w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7849w8126w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7849w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7857w8134w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7857w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8589w8866w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8589w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8672w8949w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8672w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8680w8957w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8680w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8688w8965w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8688w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8696w8973w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8696w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8704w8981w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8704w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8712w8989w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8712w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8720w8997w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8720w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8728w9005w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8728w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8736w9013w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8736w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8744w9021w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8744w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8600w8877w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8600w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8752w9029w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8752w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8760w9037w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8760w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8768w9045w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8768w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8776w9053w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8776w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8784w9061w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8784w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8792w9069w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8792w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8800w9077w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8800w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8808w9085w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8808w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8816w9093w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8816w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8824w9101w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8824w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8608w8885w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8608w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8832w9109w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8832w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8840w9117w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8840w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8848w9125w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8848w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8856w9133w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8856w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8616w8893w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8616w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8624w8901w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8624w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8632w8909w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8632w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8640w8917w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8640w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8648w8925w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8648w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8656w8933w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8656w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8664w8941w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8664w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9391w9668w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9391w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9474w9751w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9474w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9482w9759w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9482w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9490w9767w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9490w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9498w9775w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9498w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9506w9783w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9506w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9514w9791w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9514w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9522w9799w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9522w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9530w9807w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9530w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9538w9815w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9538w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9546w9823w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9546w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9402w9679w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9402w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9554w9831w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9554w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9562w9839w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9562w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9570w9847w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9570w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9578w9855w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9578w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9586w9863w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9586w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9594w9871w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9594w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9602w9879w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9602w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9610w9887w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9610w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9618w9895w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9618w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9626w9903w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9626w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9410w9687w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9410w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9634w9911w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9634w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9642w9919w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9642w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9650w9927w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9650w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9658w9935w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9658w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9418w9695w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9418w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9426w9703w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9426w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9434w9711w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9434w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9442w9719w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9442w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9450w9727w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9450w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9458w9735w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9458w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9466w9743w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9466w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10188w10465w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10188w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10271w10548w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10271w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10279w10556w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10279w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10287w10564w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10287w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10295w10572w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10295w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10303w10580w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10303w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10311w10588w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10311w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10319w10596w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10319w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10327w10604w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10327w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10335w10612w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10335w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10343w10620w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10343w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10199w10476w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10199w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10351w10628w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10351w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10359w10636w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10359w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10367w10644w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10367w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10375w10652w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10375w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10383w10660w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10383w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10391w10668w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10391w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10399w10676w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10399w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10407w10684w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10407w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10415w10692w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10415w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10423w10700w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10423w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10207w10484w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10207w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10431w10708w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10431w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10439w10716w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10439w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10447w10724w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10447w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10455w10732w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10455w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10215w10492w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10215w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10223w10500w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10223w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10231w10508w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10231w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10239w10516w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10239w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10247w10524w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10247w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10255w10532w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10255w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10263w10540w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10263w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1146w1423w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1146w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1229w1506w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1229w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1237w1514w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1237w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1245w1522w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1245w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1253w1530w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1253w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1261w1538w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1261w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1269w1546w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1269w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1277w1554w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1277w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1285w1562w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1285w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1293w1570w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1293w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1301w1578w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1301w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1157w1434w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1157w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1309w1586w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1309w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1317w1594w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1317w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1325w1602w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1325w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1333w1610w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1333w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1341w1618w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1341w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1349w1626w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1349w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1357w1634w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1357w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1365w1642w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1365w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1373w1650w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1373w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1381w1658w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1381w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1165w1442w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1165w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1389w1666w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1389w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1397w1674w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1397w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1405w1682w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1405w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1413w1690w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1413w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1173w1450w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1173w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1181w1458w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1181w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1189w1466w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1189w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1197w1474w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1197w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1205w1482w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1205w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1213w1490w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1213w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1221w1498w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1221w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1993w2270w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1993w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2076w2353w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2076w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2084w2361w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2084w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2092w2369w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2092w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2100w2377w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2100w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2108w2385w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2108w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2116w2393w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2116w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2124w2401w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2124w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2132w2409w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2132w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2140w2417w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2140w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2148w2425w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2148w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2004w2281w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2004w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2156w2433w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2156w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2164w2441w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2164w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2172w2449w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2172w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2180w2457w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2180w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2188w2465w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2188w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2196w2473w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2196w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2204w2481w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2204w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2212w2489w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2212w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2220w2497w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2220w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2228w2505w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2228w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2012w2289w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2012w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2236w2513w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2236w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2244w2521w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2244w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2252w2529w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2252w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2260w2537w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2260w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2020w2297w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2020w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2028w2305w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2028w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2036w2313w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2036w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2044w2321w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2044w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2052w2329w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2052w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2060w2337w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2060w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2068w2345w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2068w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2835w3112w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2835w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2918w3195w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2918w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2926w3203w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2926w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2934w3211w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2934w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2942w3219w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2942w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2950w3227w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2950w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2958w3235w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2958w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2966w3243w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2966w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2974w3251w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2974w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2982w3259w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2982w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2990w3267w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2990w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2846w3123w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2846w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2998w3275w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2998w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3006w3283w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3006w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3014w3291w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3014w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3022w3299w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3022w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3030w3307w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3030w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3038w3315w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3038w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3046w3323w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3046w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3054w3331w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3054w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3062w3339w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3062w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3070w3347w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3070w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2854w3131w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2854w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3078w3355w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3078w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3086w3363w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3086w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3094w3371w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3094w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3102w3379w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3102w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2862w3139w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2862w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2870w3147w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2870w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2878w3155w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2878w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2886w3163w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2886w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2894w3171w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2894w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2902w3179w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2902w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2910w3187w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2910w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3672w3949w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3672w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3755w4032w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3755w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3763w4040w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3763w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3771w4048w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3771w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3779w4056w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3779w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3787w4064w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3787w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3795w4072w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3795w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3803w4080w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3803w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3811w4088w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3811w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3819w4096w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3819w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3827w4104w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3827w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3683w3960w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3683w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3835w4112w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3835w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3843w4120w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3843w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3851w4128w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3851w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3859w4136w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3859w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3867w4144w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3867w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3875w4152w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3875w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3883w4160w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3883w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3891w4168w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3891w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3899w4176w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3899w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3907w4184w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3907w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3691w3968w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3691w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3915w4192w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3915w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3923w4200w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3923w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3931w4208w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3931w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3939w4216w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3939w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3699w3976w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3699w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3707w3984w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3707w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3715w3992w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3715w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3723w4000w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3723w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3731w4008w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3731w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3739w4016w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3739w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3747w4024w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3747w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4504w4781w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4504w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4587w4864w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4587w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4595w4872w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4595w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4603w4880w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4603w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4611w4888w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4611w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4619w4896w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4619w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4627w4904w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4627w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4635w4912w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4635w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4643w4920w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4643w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4651w4928w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4651w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4659w4936w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4659w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4515w4792w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4515w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4667w4944w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4667w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4675w4952w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4675w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4683w4960w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4683w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4691w4968w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4691w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4699w4976w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4699w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4707w4984w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4707w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4715w4992w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4715w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4723w5000w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4723w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4731w5008w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4731w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4739w5016w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4739w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4523w4800w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4523w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4747w5024w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4747w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4755w5032w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4755w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4763w5040w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4763w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4771w5048w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4771w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4531w4808w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4531w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4539w4816w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4539w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4547w4824w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4547w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4555w4832w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4555w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4563w4840w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4563w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4571w4848w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4571w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4579w4856w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4579w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5331w5608w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5331w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5414w5691w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5414w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5422w5699w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5422w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5430w5707w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5430w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5438w5715w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5438w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5446w5723w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5446w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5454w5731w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5454w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5462w5739w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5462w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5470w5747w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5470w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5478w5755w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5478w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5486w5763w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5486w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5342w5619w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5342w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5494w5771w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5494w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5502w5779w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5502w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5510w5787w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5510w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5518w5795w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5518w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5526w5803w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5526w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5534w5811w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5534w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5542w5819w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5542w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5550w5827w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5550w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5558w5835w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5558w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5566w5843w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5566w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5350w5627w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5350w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5574w5851w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5574w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5582w5859w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5582w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5590w5867w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5590w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5598w5875w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5598w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5358w5635w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5358w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5366w5643w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5366w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5374w5651w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5374w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5382w5659w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5382w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5390w5667w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5390w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5398w5675w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5398w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5406w5683w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5406w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6153w6430w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6153w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6236w6513w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6236w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6244w6521w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6244w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6252w6529w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6252w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6260w6537w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6260w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6268w6545w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6268w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6276w6553w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6276w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6284w6561w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6284w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6292w6569w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6292w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6300w6577w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6300w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6308w6585w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6308w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6164w6441w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6164w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6316w6593w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6316w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6324w6601w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6324w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6332w6609w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6332w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6340w6617w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6340w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6348w6625w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6348w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6356w6633w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6356w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6364w6641w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6364w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6372w6649w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6372w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6380w6657w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6380w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6388w6665w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6388w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6172w6449w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6172w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6396w6673w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6396w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6404w6681w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6404w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6412w6689w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6412w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6420w6697w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6420w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6180w6457w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6180w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6188w6465w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6188w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6196w6473w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6196w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6204w6481w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6204w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6212w6489w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6212w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6220w6497w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6220w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6228w6505w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6228w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6970w7247w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6970w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7053w7330w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7053w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7061w7338w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7061w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7069w7346w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7069w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7077w7354w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7077w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7085w7362w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7085w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7093w7370w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7093w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7101w7378w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7101w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7109w7386w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7109w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7117w7394w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7117w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7125w7402w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7125w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6981w7258w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6981w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7133w7410w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7133w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7141w7418w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7141w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7149w7426w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7149w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7157w7434w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7157w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7165w7442w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7165w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7173w7450w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7173w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7181w7458w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7181w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7189w7466w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7189w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7197w7474w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7197w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7205w7482w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7205w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6989w7266w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6989w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7213w7490w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7213w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7221w7498w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7221w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7229w7506w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7229w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7237w7514w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7237w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6997w7274w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6997w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7005w7282w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7005w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7013w7290w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7013w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7021w7298w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7021w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7029w7306w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7029w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7037w7314w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7037w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7045w7322w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7045w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7788w8062w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7788w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7869w8144w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7869w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7877w8152w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7877w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7885w8160w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7885w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7893w8168w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7893w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7901w8176w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7901w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7909w8184w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7909w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7917w8192w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7917w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7925w8200w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7925w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7933w8208w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7933w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7941w8216w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7941w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7797w8072w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7797w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7949w8224w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7949w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7957w8232w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7957w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7965w8240w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7965w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7973w8248w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7973w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7981w8256w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7981w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7989w8264w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7989w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7997w8272w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7997w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8005w8280w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range8005w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8013w8288w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range8013w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8021w8296w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range8021w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7805w8080w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7805w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8029w8304w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range8029w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8037w8312w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range8037w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8045w8320w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range8045w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8053w8328w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range8053w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7813w8088w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7813w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7821w8096w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7821w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7829w8104w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7829w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7837w8112w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7837w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7845w8120w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7845w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7853w8128w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7853w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7861w8136w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7861w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8595w8869w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8595w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8676w8951w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8676w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8684w8959w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8684w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8692w8967w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8692w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8700w8975w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8700w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8708w8983w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8708w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8716w8991w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8716w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8724w8999w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8724w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8732w9007w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8732w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8740w9015w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8740w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8748w9023w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8748w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8604w8879w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8604w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8756w9031w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8756w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8764w9039w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8764w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8772w9047w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8772w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8780w9055w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8780w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8788w9063w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8788w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8796w9071w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8796w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8804w9079w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8804w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8812w9087w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8812w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8820w9095w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8820w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8828w9103w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8828w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8612w8887w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8612w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8836w9111w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8836w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8844w9119w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8844w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8852w9127w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8852w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8860w9135w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8860w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8620w8895w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8620w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8628w8903w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8628w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8636w8911w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8636w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8644w8919w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8644w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8652w8927w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8652w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8660w8935w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8660w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8668w8943w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8668w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9397w9671w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9397w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9478w9753w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9478w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9486w9761w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9486w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9494w9769w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9494w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9502w9777w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9502w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9510w9785w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9510w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9518w9793w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9518w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9526w9801w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9526w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9534w9809w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9534w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9542w9817w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9542w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9550w9825w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9550w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9406w9681w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9406w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9558w9833w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9558w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9566w9841w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9566w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9574w9849w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9574w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9582w9857w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9582w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9590w9865w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9590w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9598w9873w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9598w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9606w9881w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9606w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9614w9889w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9614w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9622w9897w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9622w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9630w9905w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9630w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9414w9689w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9414w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9638w9913w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9638w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9646w9921w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9646w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9654w9929w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9654w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9662w9937w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9662w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9422w9697w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9422w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9430w9705w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9430w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9438w9713w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9438w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9446w9721w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9446w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9454w9729w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9454w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9462w9737w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9462w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9470w9745w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9470w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10194w10468w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10194w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10275w10550w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10275w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10283w10558w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10283w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10291w10566w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10291w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10299w10574w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10299w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10307w10582w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10307w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10315w10590w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10315w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10323w10598w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10323w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10331w10606w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10331w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10339w10614w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10339w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10347w10622w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10347w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10203w10478w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10203w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10355w10630w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10355w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10363w10638w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10363w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10371w10646w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10371w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10379w10654w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10379w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10387w10662w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10387w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10395w10670w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10395w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10403w10678w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10403w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10411w10686w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10411w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10419w10694w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10419w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10427w10702w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10427w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10211w10486w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10211w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10435w10710w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10435w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10443w10718w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10443w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10451w10726w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10451w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10459w10734w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10459w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10219w10494w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10219w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10227w10502w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10227w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10235w10510w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10235w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10243w10518w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10243w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10251w10526w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10251w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10259w10534w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10259w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10267w10542w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10267w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1152w1426w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1152w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1233w1508w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1233w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1241w1516w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1241w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1249w1524w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1249w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1257w1532w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1257w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1265w1540w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1265w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1273w1548w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1273w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1281w1556w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1281w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1289w1564w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1289w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1297w1572w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1297w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1305w1580w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1305w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1161w1436w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1161w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1313w1588w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1313w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1321w1596w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1321w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1329w1604w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1329w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1337w1612w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1337w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1345w1620w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1345w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1353w1628w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1353w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1361w1636w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1361w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1369w1644w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1369w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1377w1652w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1377w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1385w1660w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1385w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1169w1444w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1169w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1393w1668w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1393w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1401w1676w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1401w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1409w1684w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1409w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1417w1692w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1417w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1177w1452w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1177w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1185w1460w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1185w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1193w1468w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1193w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1201w1476w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1201w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1209w1484w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1209w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1217w1492w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1217w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1225w1500w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1225w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1999w2273w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1999w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2080w2355w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2080w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2088w2363w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2088w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2096w2371w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2096w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2104w2379w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2104w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2112w2387w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2112w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2120w2395w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2120w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2128w2403w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2128w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2136w2411w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2136w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2144w2419w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2144w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2152w2427w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2152w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2008w2283w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2008w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2160w2435w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2160w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2168w2443w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2168w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2176w2451w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2176w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2184w2459w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2184w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2192w2467w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2192w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2200w2475w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2200w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2208w2483w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2208w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2216w2491w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2216w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2224w2499w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2224w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2232w2507w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2232w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2016w2291w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2016w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2240w2515w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2240w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2248w2523w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2248w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2256w2531w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2256w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2264w2539w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2264w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2024w2299w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2024w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2032w2307w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2032w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2040w2315w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2040w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2048w2323w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2048w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2056w2331w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2056w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2064w2339w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2064w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2072w2347w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2072w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2841w3115w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2841w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2922w3197w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2922w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2930w3205w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2930w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2938w3213w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2938w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2946w3221w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2946w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2954w3229w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2954w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2962w3237w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2962w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2970w3245w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2970w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2978w3253w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2978w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2986w3261w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2986w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2994w3269w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2994w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2850w3125w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2850w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3002w3277w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3002w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3010w3285w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3010w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3018w3293w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3018w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3026w3301w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3026w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3034w3309w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3034w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3042w3317w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3042w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3050w3325w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3050w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3058w3333w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3058w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3066w3341w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3066w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3074w3349w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3074w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2858w3133w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2858w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3082w3357w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3082w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3090w3365w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3090w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3098w3373w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3098w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3106w3381w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3106w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2866w3141w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2866w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2874w3149w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2874w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2882w3157w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2882w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2890w3165w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2890w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2898w3173w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2898w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2906w3181w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2906w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2914w3189w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2914w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3678w3952w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3678w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3759w4034w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3759w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3767w4042w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3767w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3775w4050w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3775w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3783w4058w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3783w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3791w4066w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3791w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3799w4074w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3799w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3807w4082w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3807w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3815w4090w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3815w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3823w4098w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3823w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3831w4106w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3831w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3687w3962w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3687w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3839w4114w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3839w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3847w4122w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3847w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3855w4130w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3855w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3863w4138w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3863w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3871w4146w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3871w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3879w4154w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3879w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3887w4162w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3887w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3895w4170w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3895w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3903w4178w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3903w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3911w4186w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3911w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3695w3970w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3695w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3919w4194w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3919w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3927w4202w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3927w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3935w4210w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3935w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3943w4218w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3943w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3703w3978w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3703w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3711w3986w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3711w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3719w3994w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3719w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3727w4002w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3727w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3735w4010w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3735w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3743w4018w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3743w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3751w4026w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3751w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4510w4784w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4510w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4591w4866w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4591w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4599w4874w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4599w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4607w4882w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4607w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4615w4890w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4615w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4623w4898w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4623w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4631w4906w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4631w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4639w4914w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4639w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4647w4922w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4647w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4655w4930w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4655w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4663w4938w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4663w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4519w4794w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4519w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4671w4946w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4671w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4679w4954w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4679w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4687w4962w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4687w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4695w4970w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4695w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4703w4978w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4703w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4711w4986w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4711w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4719w4994w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4719w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4727w5002w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4727w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4735w5010w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4735w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4743w5018w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4743w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4527w4802w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4527w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4751w5026w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4751w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4759w5034w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4759w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4767w5042w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4767w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4775w5050w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4775w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4535w4810w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4535w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4543w4818w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4543w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4551w4826w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4551w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4559w4834w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4559w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4567w4842w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4567w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4575w4850w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4575w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4583w4858w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4583w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5337w5611w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5337w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5418w5693w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5418w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5426w5701w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5426w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5434w5709w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5434w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5442w5717w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5442w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5450w5725w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5450w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5458w5733w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5458w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5466w5741w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5466w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5474w5749w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5474w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5482w5757w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5482w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5490w5765w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5490w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5346w5621w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5346w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5498w5773w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5498w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5506w5781w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5506w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5514w5789w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5514w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5522w5797w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5522w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5530w5805w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5530w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5538w5813w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5538w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5546w5821w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5546w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5554w5829w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5554w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5562w5837w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5562w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5570w5845w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5570w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5354w5629w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5354w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5578w5853w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5578w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5586w5861w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5586w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5594w5869w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5594w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5602w5877w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5602w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5362w5637w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5362w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5370w5645w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5370w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5378w5653w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5378w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5386w5661w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5386w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5394w5669w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5394w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5402w5677w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5402w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5410w5685w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5410w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6159w6433w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6159w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6240w6515w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6240w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6248w6523w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6248w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6256w6531w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6256w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6264w6539w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6264w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6272w6547w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6272w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6280w6555w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6280w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6288w6563w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6288w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6296w6571w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6296w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6304w6579w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6304w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6312w6587w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6312w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6168w6443w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6168w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6320w6595w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6320w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6328w6603w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6328w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6336w6611w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6336w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6344w6619w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6344w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6352w6627w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6352w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6360w6635w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6360w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6368w6643w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6368w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6376w6651w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6376w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6384w6659w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6384w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6392w6667w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6392w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6176w6451w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6176w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6400w6675w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6400w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6408w6683w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6408w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6416w6691w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6416w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6424w6699w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6424w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6184w6459w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6184w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6192w6467w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6192w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6200w6475w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6200w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6208w6483w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6208w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6216w6491w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6216w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6224w6499w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6224w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6232w6507w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6232w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6976w7250w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6976w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7057w7332w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7057w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7065w7340w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7065w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7073w7348w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7073w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7081w7356w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7081w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7089w7364w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7089w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7097w7372w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7097w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7105w7380w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7105w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7113w7388w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7113w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7121w7396w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7121w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7129w7404w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7129w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6985w7260w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6985w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7137w7412w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7137w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7145w7420w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7145w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7153w7428w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7153w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7161w7436w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7161w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7169w7444w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7169w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7177w7452w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7177w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7185w7460w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7185w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7193w7468w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7193w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7201w7476w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7201w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7209w7484w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7209w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6993w7268w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6993w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7217w7492w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7217w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7225w7500w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7225w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7233w7508w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7233w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7241w7516w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7241w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7001w7276w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7001w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7009w7284w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7009w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7017w7292w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7017w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7025w7300w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7025w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7033w7308w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7033w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7041w7316w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7041w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7049w7324w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7049w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	atannode_0_w <= wire_cata_0_cordic_atan_arctan;
	atannode_10_w <= wire_cata_10_cordic_atan_arctan;
	atannode_11_w <= wire_cata_11_cordic_atan_arctan;
	atannode_12_w <= wire_cata_12_cordic_atan_arctan;
	atannode_1_w <= wire_cata_1_cordic_atan_arctan;
	atannode_2_w <= wire_cata_2_cordic_atan_arctan;
	atannode_3_w <= wire_cata_3_cordic_atan_arctan;
	atannode_4_w <= wire_cata_4_cordic_atan_arctan;
	atannode_5_w <= wire_cata_5_cordic_atan_arctan;
	atannode_6_w <= wire_cata_6_cordic_atan_arctan;
	atannode_7_w <= wire_cata_7_cordic_atan_arctan;
	atannode_8_w <= wire_cata_8_cordic_atan_arctan;
	atannode_9_w <= wire_cata_9_cordic_atan_arctan;
	delay_input_w <= (wire_x_pipeff_13_w_lg_q10744w OR wire_y_pipeff_13_w_lg_q10743w);
	delay_pipe_w <= cdaff_2;
	estimate_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10909w10918w10919w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10904w10915w10916w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10899w10912w10913w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10894w10907w10908w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10889w10902w10903w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10884w10897w10898w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10879w10892w10893w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10874w10887w10888w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10869w10882w10883w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10864w10877w10878w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10859w10872w10873w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10854w10867w10868w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10849w10862w10863w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10844w10857w10858w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10839w10852w10853w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10834w10847w10848w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10829w10842w10843w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10824w10837w10838w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10819w10832w10833w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10814w10827w10828w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10809w10822w10823w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10804w10817w10818w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10799w10812w10813w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10794w10807w10808w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10789w10802w10803w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10784w10797w10798w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10779w10792w10793w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10774w10787w10788w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10769w10782w10783w
 & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10764w10777w10778w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10758w10772w10773w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10750w10767w10768w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10759w10762w10763w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10751w10755w10756w);
	indexpointnum_w <= (OTHERS => '0');
	multiplier_input_w <= (wire_x_pipeff_13_w_lg_q10741w OR wire_y_pipeff_13_w_lg_q10740w);
	multipliernode_w <= wire_cmx_result;
	post_estimate_w <= wire_ccc_cordic_m_w_lg_estimate_w10920w;
	pre_estimate_w <= multipliernode_w(65 DOWNTO 32);
	radians_load_node_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_radians_range573w576w577w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range568w571w572w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range563w566w567w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range558w561w562w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range553w556w557w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range548w551w552w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range543w546w547w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range538w541w542w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range533w536w537w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range528w531w532w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range523w526w527w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range518w521w522w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range513w516w517w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range508w511w512w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range503w506w507w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range498w501w502w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range493w496w497w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range488w491w492w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range483w486w487w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range478w481w482w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range473w476w477w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range468w471w472w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range463w466w467w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range458w461w462w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range453w456w457w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range448w451w452w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range443w446w447w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range438w441w442w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range433w436w437w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range428w431w432w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range423w426w427w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range418w421w422w & wire_ccc_cordic_m_w_lg_w_radians_range415w417w & wire_ccc_cordic_m_w_lg_w_radians_range410w413w);
	sincos <= sincosff;
	startindex_w <= wire_ccc_cordic_m_w_lg_indexpointnum_w409w;
	x_pipenode_10_w <= wire_x_pipenode_10_add_result;
	x_pipenode_11_w <= wire_x_pipenode_11_add_result;
	x_pipenode_12_w <= wire_x_pipenode_12_add_result;
	x_pipenode_13_w <= wire_x_pipenode_13_add_result;
	x_pipenode_2_w <= wire_x_pipenode_2_add_result;
	x_pipenode_3_w <= wire_x_pipenode_3_add_result;
	x_pipenode_4_w <= wire_x_pipenode_4_add_result;
	x_pipenode_5_w <= wire_x_pipenode_5_add_result;
	x_pipenode_6_w <= wire_x_pipenode_6_add_result;
	x_pipenode_7_w <= wire_x_pipenode_7_add_result;
	x_pipenode_8_w <= wire_x_pipenode_8_add_result;
	x_pipenode_9_w <= wire_x_pipenode_9_add_result;
	x_prenode_10_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7542w8051w8052w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7540w8043w8044w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7538w8035w8036w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7536w8027w8028w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7534w8019w8020w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7532w8011w8012w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7530w8003w8004w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7528w7995w7996w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7522w7987w7988w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7711w7979w7980w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7706w7971w7972w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7700w7963w7964w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7694w7955w7956w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7688w7947w7948w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7682w7939w7940w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7676w7931w7932w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7670w7923w7924w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7664w7915w7916w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7658w7907w7908w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7652w7899w7900w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7646w7891w7892w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7640w7883w7884w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7634w7875w7876w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7628w7867w7868w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7622w7859w7860w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7616w7851w7852w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7610w7843w7844w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7604w7835w7836w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7598w7827w7828w
 & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7592w7819w7820w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7586w7811w7812w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7580w7803w7804w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7574w7795w7796w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7569w7785w7786w);
	x_prenode_11_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8356w8858w8859w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8354w8850w8851w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8352w8842w8843w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8350w8834w8835w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8348w8826w8827w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8346w8818w8819w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8344w8810w8811w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8342w8802w8803w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8340w8794w8795w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8334w8786w8787w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8521w8778w8779w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8516w8770w8771w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8510w8762w8763w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8504w8754w8755w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8498w8746w8747w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8492w8738w8739w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8486w8730w8731w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8480w8722w8723w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8474w8714w8715w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8468w8706w8707w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8462w8698w8699w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8456w8690w8691w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8450w8682w8683w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8444w8674w8675w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8438w8666w8667w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8432w8658w8659w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8426w8650w8651w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8420w8642w8643w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8414w8634w8635w
 & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8408w8626w8627w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8402w8618w8619w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8396w8610w8611w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8390w8602w8603w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8385w8592w8593w);
	x_prenode_12_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9165w9660w9661w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9163w9652w9653w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9161w9644w9645w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9159w9636w9637w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9157w9628w9629w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9155w9620w9621w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9153w9612w9613w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9151w9604w9605w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9149w9596w9597w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9147w9588w9589w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9141w9580w9581w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9326w9572w9573w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9321w9564w9565w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9315w9556w9557w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9309w9548w9549w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9303w9540w9541w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9297w9532w9533w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9291w9524w9525w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9285w9516w9517w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9279w9508w9509w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9273w9500w9501w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9267w9492w9493w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9261w9484w9485w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9255w9476w9477w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9249w9468w9469w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9243w9460w9461w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9237w9452w9453w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9231w9444w9445w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9225w9436w9437w
 & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9219w9428w9429w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9213w9420w9421w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9207w9412w9413w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9201w9404w9405w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9196w9394w9395w);
	x_prenode_13_w <= ( wire_ccc_cordic_m_w10458w & wire_ccc_cordic_m_w10450w & wire_ccc_cordic_m_w10442w & wire_ccc_cordic_m_w10434w & wire_ccc_cordic_m_w10426w & wire_ccc_cordic_m_w10418w & wire_ccc_cordic_m_w10410w & wire_ccc_cordic_m_w10402w & wire_ccc_cordic_m_w10394w & wire_ccc_cordic_m_w10386w & wire_ccc_cordic_m_w10378w & wire_ccc_cordic_m_w10370w & wire_ccc_cordic_m_w10362w & wire_ccc_cordic_m_w10354w & wire_ccc_cordic_m_w10346w & wire_ccc_cordic_m_w10338w & wire_ccc_cordic_m_w10330w & wire_ccc_cordic_m_w10322w & wire_ccc_cordic_m_w10314w & wire_ccc_cordic_m_w10306w & wire_ccc_cordic_m_w10298w & wire_ccc_cordic_m_w10290w & wire_ccc_cordic_m_w10282w & wire_ccc_cordic_m_w10274w & wire_ccc_cordic_m_w10266w & wire_ccc_cordic_m_w10258w & wire_ccc_cordic_m_w10250w & wire_ccc_cordic_m_w10242w & wire_ccc_cordic_m_w10234w & wire_ccc_cordic_m_w10226w & wire_ccc_cordic_m_w10218w & wire_ccc_cordic_m_w10210w & wire_ccc_cordic_m_w10202w & wire_ccc_cordic_m_w10192w);
	x_prenode_2_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range846w1415w1416w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1051w1407w1408w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1046w1399w1400w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1040w1391w1392w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1034w1383w1384w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1028w1375w1376w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1022w1367w1368w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1016w1359w1360w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1010w1351w1352w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1004w1343w1344w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range998w1335w1336w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range992w1327w1328w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range986w1319w1320w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range980w1311w1312w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range974w1303w1304w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range968w1295w1296w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range962w1287w1288w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range956w1279w1280w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range950w1271w1272w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range944w1263w1264w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range938w1255w1256w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range932w1247w1248w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range926w1239w1240w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range920w1231w1232w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range914w1223w1224w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range908w1215w1216w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range902w1207w1208w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range896w1199w1200w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range890w1191w1192w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range884w1183w1184w
 & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range878w1175w1176w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range872w1167w1168w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range866w1159w1160w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range861w1149w1150w);
	x_prenode_3_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1704w2262w2263w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1698w2254w2255w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1901w2246w2247w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1896w2238w2239w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1890w2230w2231w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1884w2222w2223w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1878w2214w2215w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1872w2206w2207w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1866w2198w2199w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1860w2190w2191w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1854w2182w2183w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1848w2174w2175w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1842w2166w2167w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1836w2158w2159w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1830w2150w2151w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1824w2142w2143w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1818w2134w2135w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1812w2126w2127w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1806w2118w2119w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1800w2110w2111w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1794w2102w2103w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1788w2094w2095w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1782w2086w2087w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1776w2078w2079w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1770w2070w2071w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1764w2062w2063w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1758w2054w2055w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1752w2046w2047w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1746w2038w2039w 
& wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1740w2030w2031w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1734w2022w2023w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1728w2014w2015w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1722w2006w2007w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1717w1996w1997w);
	x_prenode_4_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2553w3104w3105w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2551w3096w3097w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2545w3088w3089w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2746w3080w3081w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2741w3072w3073w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2735w3064w3065w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2729w3056w3057w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2723w3048w3049w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2717w3040w3041w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2711w3032w3033w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2705w3024w3025w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2699w3016w3017w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2693w3008w3009w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2687w3000w3001w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2681w2992w2993w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2675w2984w2985w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2669w2976w2977w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2663w2968w2969w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2657w2960w2961w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2651w2952w2953w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2645w2944w2945w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2639w2936w2937w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2633w2928w2929w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2627w2920w2921w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2621w2912w2913w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2615w2904w2905w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2609w2896w2897w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2603w2888w2889w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2597w2880w2881w 
& wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2591w2872w2873w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2585w2864w2865w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2579w2856w2857w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2573w2848w2849w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2568w2838w2839w);
	x_prenode_5_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3397w3941w3942w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3395w3933w3934w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3393w3925w3926w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3387w3917w3918w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3586w3909w3910w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3581w3901w3902w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3575w3893w3894w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3569w3885w3886w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3563w3877w3878w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3557w3869w3870w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3551w3861w3862w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3545w3853w3854w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3539w3845w3846w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3533w3837w3838w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3527w3829w3830w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3521w3821w3822w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3515w3813w3814w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3509w3805w3806w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3503w3797w3798w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3497w3789w3790w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3491w3781w3782w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3485w3773w3774w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3479w3765w3766w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3473w3757w3758w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3467w3749w3750w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3461w3741w3742w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3455w3733w3734w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3449w3725w3726w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3443w3717w3718w 
& wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3437w3709w3710w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3431w3701w3702w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3425w3693w3694w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3419w3685w3686w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3414w3675w3676w);
	x_prenode_6_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4236w4773w4774w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4234w4765w4766w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4232w4757w4758w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4230w4749w4750w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4224w4741w4742w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4421w4733w4734w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4416w4725w4726w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4410w4717w4718w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4404w4709w4710w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4398w4701w4702w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4392w4693w4694w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4386w4685w4686w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4380w4677w4678w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4374w4669w4670w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4368w4661w4662w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4362w4653w4654w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4356w4645w4646w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4350w4637w4638w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4344w4629w4630w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4338w4621w4622w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4332w4613w4614w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4326w4605w4606w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4320w4597w4598w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4314w4589w4590w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4308w4581w4582w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4302w4573w4574w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4296w4565w4566w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4290w4557w4558w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4284w4549w4550w 
& wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4278w4541w4542w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4272w4533w4534w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4266w4525w4526w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4260w4517w4518w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4255w4507w4508w);
	x_prenode_7_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5070w5600w5601w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5068w5592w5593w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5066w5584w5585w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5064w5576w5577w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5062w5568w5569w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5056w5560w5561w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5251w5552w5553w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5246w5544w5545w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5240w5536w5537w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5234w5528w5529w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5228w5520w5521w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5222w5512w5513w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5216w5504w5505w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5210w5496w5497w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5204w5488w5489w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5198w5480w5481w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5192w5472w5473w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5186w5464w5465w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5180w5456w5457w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5174w5448w5449w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5168w5440w5441w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5162w5432w5433w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5156w5424w5425w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5150w5416w5417w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5144w5408w5409w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5138w5400w5401w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5132w5392w5393w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5126w5384w5385w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5120w5376w5377w 
& wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5114w5368w5369w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5108w5360w5361w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5102w5352w5353w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5096w5344w5345w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5091w5334w5335w);
	x_prenode_8_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5899w6422w6423w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5897w6414w6415w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5895w6406w6407w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5893w6398w6399w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5891w6390w6391w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5889w6382w6383w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5883w6374w6375w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6076w6366w6367w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6071w6358w6359w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6065w6350w6351w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6059w6342w6343w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6053w6334w6335w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6047w6326w6327w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6041w6318w6319w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6035w6310w6311w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6029w6302w6303w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6023w6294w6295w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6017w6286w6287w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6011w6278w6279w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6005w6270w6271w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5999w6262w6263w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5993w6254w6255w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5987w6246w6247w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5981w6238w6239w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5975w6230w6231w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5969w6222w6223w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5963w6214w6215w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5957w6206w6207w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5951w6198w6199w 
& wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5945w6190w6191w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5939w6182w6183w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5933w6174w6175w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5927w6166w6167w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5922w6156w6157w);
	x_prenode_9_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6723w7239w7240w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6721w7231w7232w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6719w7223w7224w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6717w7215w7216w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6715w7207w7208w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6713w7199w7200w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6711w7191w7192w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6705w7183w7184w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6896w7175w7176w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6891w7167w7168w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6885w7159w7160w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6879w7151w7152w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6873w7143w7144w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6867w7135w7136w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6861w7127w7128w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6855w7119w7120w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6849w7111w7112w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6843w7103w7104w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6837w7095w7096w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6831w7087w7088w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6825w7079w7080w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6819w7071w7072w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6813w7063w7064w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6807w7055w7056w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6801w7047w7048w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6795w7039w7040w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6789w7031w7032w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6783w7023w7024w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6777w7015w7016w 
& wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6771w7007w7008w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6765w6999w7000w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6759w6991w6992w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6753w6983w6984w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6748w6973w6974w);
	x_prenodeone_10_w <= ( wire_y_pipeff_9_w_lg_w_q_range7521w7523w & wire_y_pipeff_9_w_lg_w_q_range7521w7523w & wire_y_pipeff_9_w_lg_w_q_range7521w7523w & wire_y_pipeff_9_w_lg_w_q_range7521w7523w & wire_y_pipeff_9_w_lg_w_q_range7521w7523w & wire_y_pipeff_9_w_lg_w_q_range7521w7523w & wire_y_pipeff_9_w_lg_w_q_range7521w7523w & wire_y_pipeff_9_w_lg_w_q_range7521w7523w & wire_y_pipeff_9_w_lg_w_q_range7521w7523w & wire_y_pipeff_9_w_lg_w_q_range7521w7523w & wire_y_pipeff_9_w_lg_w_q_range7705w7707w & wire_y_pipeff_9_w_lg_w_q_range7699w7701w & wire_y_pipeff_9_w_lg_w_q_range7693w7695w & wire_y_pipeff_9_w_lg_w_q_range7687w7689w & wire_y_pipeff_9_w_lg_w_q_range7681w7683w & wire_y_pipeff_9_w_lg_w_q_range7675w7677w & wire_y_pipeff_9_w_lg_w_q_range7669w7671w & wire_y_pipeff_9_w_lg_w_q_range7663w7665w & wire_y_pipeff_9_w_lg_w_q_range7657w7659w & wire_y_pipeff_9_w_lg_w_q_range7651w7653w & wire_y_pipeff_9_w_lg_w_q_range7645w7647w & wire_y_pipeff_9_w_lg_w_q_range7639w7641w & wire_y_pipeff_9_w_lg_w_q_range7633w7635w & wire_y_pipeff_9_w_lg_w_q_range7627w7629w & wire_y_pipeff_9_w_lg_w_q_range7621w7623w & wire_y_pipeff_9_w_lg_w_q_range7615w7617w & wire_y_pipeff_9_w_lg_w_q_range7609w7611w & wire_y_pipeff_9_w_lg_w_q_range7603w7605w & wire_y_pipeff_9_w_lg_w_q_range7597w7599w & wire_y_pipeff_9_w_lg_w_q_range7591w7593w & wire_y_pipeff_9_w_lg_w_q_range7585w7587w & wire_y_pipeff_9_w_lg_w_q_range7579w7581w & wire_y_pipeff_9_w_lg_w_q_range7573w7575w & wire_y_pipeff_9_w_lg_w_q_range7568w7570w);
	x_prenodeone_11_w <= ( wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8515w8517w & wire_y_pipeff_10_w_lg_w_q_range8509w8511w & wire_y_pipeff_10_w_lg_w_q_range8503w8505w & wire_y_pipeff_10_w_lg_w_q_range8497w8499w & wire_y_pipeff_10_w_lg_w_q_range8491w8493w & wire_y_pipeff_10_w_lg_w_q_range8485w8487w & wire_y_pipeff_10_w_lg_w_q_range8479w8481w & wire_y_pipeff_10_w_lg_w_q_range8473w8475w & wire_y_pipeff_10_w_lg_w_q_range8467w8469w & wire_y_pipeff_10_w_lg_w_q_range8461w8463w & wire_y_pipeff_10_w_lg_w_q_range8455w8457w & wire_y_pipeff_10_w_lg_w_q_range8449w8451w & wire_y_pipeff_10_w_lg_w_q_range8443w8445w & wire_y_pipeff_10_w_lg_w_q_range8437w8439w & wire_y_pipeff_10_w_lg_w_q_range8431w8433w & wire_y_pipeff_10_w_lg_w_q_range8425w8427w & wire_y_pipeff_10_w_lg_w_q_range8419w8421w & wire_y_pipeff_10_w_lg_w_q_range8413w8415w & wire_y_pipeff_10_w_lg_w_q_range8407w8409w & wire_y_pipeff_10_w_lg_w_q_range8401w8403w & wire_y_pipeff_10_w_lg_w_q_range8395w8397w & wire_y_pipeff_10_w_lg_w_q_range8389w8391w & wire_y_pipeff_10_w_lg_w_q_range8384w8386w);
	x_prenodeone_12_w <= ( wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9320w9322w & wire_y_pipeff_11_w_lg_w_q_range9314w9316w & wire_y_pipeff_11_w_lg_w_q_range9308w9310w & wire_y_pipeff_11_w_lg_w_q_range9302w9304w & wire_y_pipeff_11_w_lg_w_q_range9296w9298w & wire_y_pipeff_11_w_lg_w_q_range9290w9292w & wire_y_pipeff_11_w_lg_w_q_range9284w9286w & wire_y_pipeff_11_w_lg_w_q_range9278w9280w & wire_y_pipeff_11_w_lg_w_q_range9272w9274w & wire_y_pipeff_11_w_lg_w_q_range9266w9268w & wire_y_pipeff_11_w_lg_w_q_range9260w9262w & wire_y_pipeff_11_w_lg_w_q_range9254w9256w & wire_y_pipeff_11_w_lg_w_q_range9248w9250w & wire_y_pipeff_11_w_lg_w_q_range9242w9244w & wire_y_pipeff_11_w_lg_w_q_range9236w9238w & wire_y_pipeff_11_w_lg_w_q_range9230w9232w & wire_y_pipeff_11_w_lg_w_q_range9224w9226w & wire_y_pipeff_11_w_lg_w_q_range9218w9220w & wire_y_pipeff_11_w_lg_w_q_range9212w9214w & wire_y_pipeff_11_w_lg_w_q_range9206w9208w & wire_y_pipeff_11_w_lg_w_q_range9200w9202w & wire_y_pipeff_11_w_lg_w_q_range9195w9197w);
	x_prenodeone_13_w <= ( wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range10120w10122w & wire_y_pipeff_12_w_lg_w_q_range10114w10116w & wire_y_pipeff_12_w_lg_w_q_range10108w10110w & wire_y_pipeff_12_w_lg_w_q_range10102w10104w & wire_y_pipeff_12_w_lg_w_q_range10096w10098w & wire_y_pipeff_12_w_lg_w_q_range10090w10092w & wire_y_pipeff_12_w_lg_w_q_range10084w10086w & wire_y_pipeff_12_w_lg_w_q_range10078w10080w & wire_y_pipeff_12_w_lg_w_q_range10072w10074w & wire_y_pipeff_12_w_lg_w_q_range10066w10068w & wire_y_pipeff_12_w_lg_w_q_range10060w10062w & wire_y_pipeff_12_w_lg_w_q_range10054w10056w & wire_y_pipeff_12_w_lg_w_q_range10048w10050w & wire_y_pipeff_12_w_lg_w_q_range10042w10044w & wire_y_pipeff_12_w_lg_w_q_range10036w10038w & wire_y_pipeff_12_w_lg_w_q_range10030w10032w & wire_y_pipeff_12_w_lg_w_q_range10024w10026w & wire_y_pipeff_12_w_lg_w_q_range10018w10020w & wire_y_pipeff_12_w_lg_w_q_range10012w10014w & wire_y_pipeff_12_w_lg_w_q_range10006w10008w & wire_y_pipeff_12_w_lg_w_q_range10001w10003w);
	x_prenodeone_2_w <= ( wire_y_pipeff_1_w_lg_w_q_range845w847w & wire_y_pipeff_1_w_lg_w_q_range845w847w & wire_y_pipeff_1_w_lg_w_q_range1045w1047w & wire_y_pipeff_1_w_lg_w_q_range1039w1041w & wire_y_pipeff_1_w_lg_w_q_range1033w1035w & wire_y_pipeff_1_w_lg_w_q_range1027w1029w & wire_y_pipeff_1_w_lg_w_q_range1021w1023w & wire_y_pipeff_1_w_lg_w_q_range1015w1017w & wire_y_pipeff_1_w_lg_w_q_range1009w1011w & wire_y_pipeff_1_w_lg_w_q_range1003w1005w & wire_y_pipeff_1_w_lg_w_q_range997w999w & wire_y_pipeff_1_w_lg_w_q_range991w993w & wire_y_pipeff_1_w_lg_w_q_range985w987w & wire_y_pipeff_1_w_lg_w_q_range979w981w & wire_y_pipeff_1_w_lg_w_q_range973w975w & wire_y_pipeff_1_w_lg_w_q_range967w969w & wire_y_pipeff_1_w_lg_w_q_range961w963w & wire_y_pipeff_1_w_lg_w_q_range955w957w & wire_y_pipeff_1_w_lg_w_q_range949w951w & wire_y_pipeff_1_w_lg_w_q_range943w945w & wire_y_pipeff_1_w_lg_w_q_range937w939w & wire_y_pipeff_1_w_lg_w_q_range931w933w & wire_y_pipeff_1_w_lg_w_q_range925w927w & wire_y_pipeff_1_w_lg_w_q_range919w921w & wire_y_pipeff_1_w_lg_w_q_range913w915w & wire_y_pipeff_1_w_lg_w_q_range907w909w & wire_y_pipeff_1_w_lg_w_q_range901w903w & wire_y_pipeff_1_w_lg_w_q_range895w897w & wire_y_pipeff_1_w_lg_w_q_range889w891w & wire_y_pipeff_1_w_lg_w_q_range883w885w & wire_y_pipeff_1_w_lg_w_q_range877w879w & wire_y_pipeff_1_w_lg_w_q_range871w873w & wire_y_pipeff_1_w_lg_w_q_range865w867w & wire_y_pipeff_1_w_lg_w_q_range860w862w);
	x_prenodeone_3_w <= ( wire_y_pipeff_2_w_lg_w_q_range1697w1699w & wire_y_pipeff_2_w_lg_w_q_range1697w1699w & wire_y_pipeff_2_w_lg_w_q_range1697w1699w & wire_y_pipeff_2_w_lg_w_q_range1895w1897w & wire_y_pipeff_2_w_lg_w_q_range1889w1891w & wire_y_pipeff_2_w_lg_w_q_range1883w1885w & wire_y_pipeff_2_w_lg_w_q_range1877w1879w & wire_y_pipeff_2_w_lg_w_q_range1871w1873w & wire_y_pipeff_2_w_lg_w_q_range1865w1867w & wire_y_pipeff_2_w_lg_w_q_range1859w1861w & wire_y_pipeff_2_w_lg_w_q_range1853w1855w & wire_y_pipeff_2_w_lg_w_q_range1847w1849w & wire_y_pipeff_2_w_lg_w_q_range1841w1843w & wire_y_pipeff_2_w_lg_w_q_range1835w1837w & wire_y_pipeff_2_w_lg_w_q_range1829w1831w & wire_y_pipeff_2_w_lg_w_q_range1823w1825w & wire_y_pipeff_2_w_lg_w_q_range1817w1819w & wire_y_pipeff_2_w_lg_w_q_range1811w1813w & wire_y_pipeff_2_w_lg_w_q_range1805w1807w & wire_y_pipeff_2_w_lg_w_q_range1799w1801w & wire_y_pipeff_2_w_lg_w_q_range1793w1795w & wire_y_pipeff_2_w_lg_w_q_range1787w1789w & wire_y_pipeff_2_w_lg_w_q_range1781w1783w & wire_y_pipeff_2_w_lg_w_q_range1775w1777w & wire_y_pipeff_2_w_lg_w_q_range1769w1771w & wire_y_pipeff_2_w_lg_w_q_range1763w1765w & wire_y_pipeff_2_w_lg_w_q_range1757w1759w & wire_y_pipeff_2_w_lg_w_q_range1751w1753w & wire_y_pipeff_2_w_lg_w_q_range1745w1747w & wire_y_pipeff_2_w_lg_w_q_range1739w1741w & wire_y_pipeff_2_w_lg_w_q_range1733w1735w & wire_y_pipeff_2_w_lg_w_q_range1727w1729w & wire_y_pipeff_2_w_lg_w_q_range1721w1723w & wire_y_pipeff_2_w_lg_w_q_range1716w1718w);
	x_prenodeone_4_w <= ( wire_y_pipeff_3_w_lg_w_q_range2544w2546w & wire_y_pipeff_3_w_lg_w_q_range2544w2546w & wire_y_pipeff_3_w_lg_w_q_range2544w2546w & wire_y_pipeff_3_w_lg_w_q_range2544w2546w & wire_y_pipeff_3_w_lg_w_q_range2740w2742w & wire_y_pipeff_3_w_lg_w_q_range2734w2736w & wire_y_pipeff_3_w_lg_w_q_range2728w2730w & wire_y_pipeff_3_w_lg_w_q_range2722w2724w & wire_y_pipeff_3_w_lg_w_q_range2716w2718w & wire_y_pipeff_3_w_lg_w_q_range2710w2712w & wire_y_pipeff_3_w_lg_w_q_range2704w2706w & wire_y_pipeff_3_w_lg_w_q_range2698w2700w & wire_y_pipeff_3_w_lg_w_q_range2692w2694w & wire_y_pipeff_3_w_lg_w_q_range2686w2688w & wire_y_pipeff_3_w_lg_w_q_range2680w2682w & wire_y_pipeff_3_w_lg_w_q_range2674w2676w & wire_y_pipeff_3_w_lg_w_q_range2668w2670w & wire_y_pipeff_3_w_lg_w_q_range2662w2664w & wire_y_pipeff_3_w_lg_w_q_range2656w2658w & wire_y_pipeff_3_w_lg_w_q_range2650w2652w & wire_y_pipeff_3_w_lg_w_q_range2644w2646w & wire_y_pipeff_3_w_lg_w_q_range2638w2640w & wire_y_pipeff_3_w_lg_w_q_range2632w2634w & wire_y_pipeff_3_w_lg_w_q_range2626w2628w & wire_y_pipeff_3_w_lg_w_q_range2620w2622w & wire_y_pipeff_3_w_lg_w_q_range2614w2616w & wire_y_pipeff_3_w_lg_w_q_range2608w2610w & wire_y_pipeff_3_w_lg_w_q_range2602w2604w & wire_y_pipeff_3_w_lg_w_q_range2596w2598w & wire_y_pipeff_3_w_lg_w_q_range2590w2592w & wire_y_pipeff_3_w_lg_w_q_range2584w2586w & wire_y_pipeff_3_w_lg_w_q_range2578w2580w & wire_y_pipeff_3_w_lg_w_q_range2572w2574w & wire_y_pipeff_3_w_lg_w_q_range2567w2569w);
	x_prenodeone_5_w <= ( wire_y_pipeff_4_w_lg_w_q_range3386w3388w & wire_y_pipeff_4_w_lg_w_q_range3386w3388w & wire_y_pipeff_4_w_lg_w_q_range3386w3388w & wire_y_pipeff_4_w_lg_w_q_range3386w3388w & wire_y_pipeff_4_w_lg_w_q_range3386w3388w & wire_y_pipeff_4_w_lg_w_q_range3580w3582w & wire_y_pipeff_4_w_lg_w_q_range3574w3576w & wire_y_pipeff_4_w_lg_w_q_range3568w3570w & wire_y_pipeff_4_w_lg_w_q_range3562w3564w & wire_y_pipeff_4_w_lg_w_q_range3556w3558w & wire_y_pipeff_4_w_lg_w_q_range3550w3552w & wire_y_pipeff_4_w_lg_w_q_range3544w3546w & wire_y_pipeff_4_w_lg_w_q_range3538w3540w & wire_y_pipeff_4_w_lg_w_q_range3532w3534w & wire_y_pipeff_4_w_lg_w_q_range3526w3528w & wire_y_pipeff_4_w_lg_w_q_range3520w3522w & wire_y_pipeff_4_w_lg_w_q_range3514w3516w & wire_y_pipeff_4_w_lg_w_q_range3508w3510w & wire_y_pipeff_4_w_lg_w_q_range3502w3504w & wire_y_pipeff_4_w_lg_w_q_range3496w3498w & wire_y_pipeff_4_w_lg_w_q_range3490w3492w & wire_y_pipeff_4_w_lg_w_q_range3484w3486w & wire_y_pipeff_4_w_lg_w_q_range3478w3480w & wire_y_pipeff_4_w_lg_w_q_range3472w3474w & wire_y_pipeff_4_w_lg_w_q_range3466w3468w & wire_y_pipeff_4_w_lg_w_q_range3460w3462w & wire_y_pipeff_4_w_lg_w_q_range3454w3456w & wire_y_pipeff_4_w_lg_w_q_range3448w3450w & wire_y_pipeff_4_w_lg_w_q_range3442w3444w & wire_y_pipeff_4_w_lg_w_q_range3436w3438w & wire_y_pipeff_4_w_lg_w_q_range3430w3432w & wire_y_pipeff_4_w_lg_w_q_range3424w3426w & wire_y_pipeff_4_w_lg_w_q_range3418w3420w & wire_y_pipeff_4_w_lg_w_q_range3413w3415w);
	x_prenodeone_6_w <= ( wire_y_pipeff_5_w_lg_w_q_range4223w4225w & wire_y_pipeff_5_w_lg_w_q_range4223w4225w & wire_y_pipeff_5_w_lg_w_q_range4223w4225w & wire_y_pipeff_5_w_lg_w_q_range4223w4225w & wire_y_pipeff_5_w_lg_w_q_range4223w4225w & wire_y_pipeff_5_w_lg_w_q_range4223w4225w & wire_y_pipeff_5_w_lg_w_q_range4415w4417w & wire_y_pipeff_5_w_lg_w_q_range4409w4411w & wire_y_pipeff_5_w_lg_w_q_range4403w4405w & wire_y_pipeff_5_w_lg_w_q_range4397w4399w & wire_y_pipeff_5_w_lg_w_q_range4391w4393w & wire_y_pipeff_5_w_lg_w_q_range4385w4387w & wire_y_pipeff_5_w_lg_w_q_range4379w4381w & wire_y_pipeff_5_w_lg_w_q_range4373w4375w & wire_y_pipeff_5_w_lg_w_q_range4367w4369w & wire_y_pipeff_5_w_lg_w_q_range4361w4363w & wire_y_pipeff_5_w_lg_w_q_range4355w4357w & wire_y_pipeff_5_w_lg_w_q_range4349w4351w & wire_y_pipeff_5_w_lg_w_q_range4343w4345w & wire_y_pipeff_5_w_lg_w_q_range4337w4339w & wire_y_pipeff_5_w_lg_w_q_range4331w4333w & wire_y_pipeff_5_w_lg_w_q_range4325w4327w & wire_y_pipeff_5_w_lg_w_q_range4319w4321w & wire_y_pipeff_5_w_lg_w_q_range4313w4315w & wire_y_pipeff_5_w_lg_w_q_range4307w4309w & wire_y_pipeff_5_w_lg_w_q_range4301w4303w & wire_y_pipeff_5_w_lg_w_q_range4295w4297w & wire_y_pipeff_5_w_lg_w_q_range4289w4291w & wire_y_pipeff_5_w_lg_w_q_range4283w4285w & wire_y_pipeff_5_w_lg_w_q_range4277w4279w & wire_y_pipeff_5_w_lg_w_q_range4271w4273w & wire_y_pipeff_5_w_lg_w_q_range4265w4267w & wire_y_pipeff_5_w_lg_w_q_range4259w4261w & wire_y_pipeff_5_w_lg_w_q_range4254w4256w);
	x_prenodeone_7_w <= ( wire_y_pipeff_6_w_lg_w_q_range5055w5057w & wire_y_pipeff_6_w_lg_w_q_range5055w5057w & wire_y_pipeff_6_w_lg_w_q_range5055w5057w & wire_y_pipeff_6_w_lg_w_q_range5055w5057w & wire_y_pipeff_6_w_lg_w_q_range5055w5057w & wire_y_pipeff_6_w_lg_w_q_range5055w5057w & wire_y_pipeff_6_w_lg_w_q_range5055w5057w & wire_y_pipeff_6_w_lg_w_q_range5245w5247w & wire_y_pipeff_6_w_lg_w_q_range5239w5241w & wire_y_pipeff_6_w_lg_w_q_range5233w5235w & wire_y_pipeff_6_w_lg_w_q_range5227w5229w & wire_y_pipeff_6_w_lg_w_q_range5221w5223w & wire_y_pipeff_6_w_lg_w_q_range5215w5217w & wire_y_pipeff_6_w_lg_w_q_range5209w5211w & wire_y_pipeff_6_w_lg_w_q_range5203w5205w & wire_y_pipeff_6_w_lg_w_q_range5197w5199w & wire_y_pipeff_6_w_lg_w_q_range5191w5193w & wire_y_pipeff_6_w_lg_w_q_range5185w5187w & wire_y_pipeff_6_w_lg_w_q_range5179w5181w & wire_y_pipeff_6_w_lg_w_q_range5173w5175w & wire_y_pipeff_6_w_lg_w_q_range5167w5169w & wire_y_pipeff_6_w_lg_w_q_range5161w5163w & wire_y_pipeff_6_w_lg_w_q_range5155w5157w & wire_y_pipeff_6_w_lg_w_q_range5149w5151w & wire_y_pipeff_6_w_lg_w_q_range5143w5145w & wire_y_pipeff_6_w_lg_w_q_range5137w5139w & wire_y_pipeff_6_w_lg_w_q_range5131w5133w & wire_y_pipeff_6_w_lg_w_q_range5125w5127w & wire_y_pipeff_6_w_lg_w_q_range5119w5121w & wire_y_pipeff_6_w_lg_w_q_range5113w5115w & wire_y_pipeff_6_w_lg_w_q_range5107w5109w & wire_y_pipeff_6_w_lg_w_q_range5101w5103w & wire_y_pipeff_6_w_lg_w_q_range5095w5097w & wire_y_pipeff_6_w_lg_w_q_range5090w5092w);
	x_prenodeone_8_w <= ( wire_y_pipeff_7_w_lg_w_q_range5882w5884w & wire_y_pipeff_7_w_lg_w_q_range5882w5884w & wire_y_pipeff_7_w_lg_w_q_range5882w5884w & wire_y_pipeff_7_w_lg_w_q_range5882w5884w & wire_y_pipeff_7_w_lg_w_q_range5882w5884w & wire_y_pipeff_7_w_lg_w_q_range5882w5884w & wire_y_pipeff_7_w_lg_w_q_range5882w5884w & wire_y_pipeff_7_w_lg_w_q_range5882w5884w & wire_y_pipeff_7_w_lg_w_q_range6070w6072w & wire_y_pipeff_7_w_lg_w_q_range6064w6066w & wire_y_pipeff_7_w_lg_w_q_range6058w6060w & wire_y_pipeff_7_w_lg_w_q_range6052w6054w & wire_y_pipeff_7_w_lg_w_q_range6046w6048w & wire_y_pipeff_7_w_lg_w_q_range6040w6042w & wire_y_pipeff_7_w_lg_w_q_range6034w6036w & wire_y_pipeff_7_w_lg_w_q_range6028w6030w & wire_y_pipeff_7_w_lg_w_q_range6022w6024w & wire_y_pipeff_7_w_lg_w_q_range6016w6018w & wire_y_pipeff_7_w_lg_w_q_range6010w6012w & wire_y_pipeff_7_w_lg_w_q_range6004w6006w & wire_y_pipeff_7_w_lg_w_q_range5998w6000w & wire_y_pipeff_7_w_lg_w_q_range5992w5994w & wire_y_pipeff_7_w_lg_w_q_range5986w5988w & wire_y_pipeff_7_w_lg_w_q_range5980w5982w & wire_y_pipeff_7_w_lg_w_q_range5974w5976w & wire_y_pipeff_7_w_lg_w_q_range5968w5970w & wire_y_pipeff_7_w_lg_w_q_range5962w5964w & wire_y_pipeff_7_w_lg_w_q_range5956w5958w & wire_y_pipeff_7_w_lg_w_q_range5950w5952w & wire_y_pipeff_7_w_lg_w_q_range5944w5946w & wire_y_pipeff_7_w_lg_w_q_range5938w5940w & wire_y_pipeff_7_w_lg_w_q_range5932w5934w & wire_y_pipeff_7_w_lg_w_q_range5926w5928w & wire_y_pipeff_7_w_lg_w_q_range5921w5923w);
	x_prenodeone_9_w <= ( wire_y_pipeff_8_w_lg_w_q_range6704w6706w & wire_y_pipeff_8_w_lg_w_q_range6704w6706w & wire_y_pipeff_8_w_lg_w_q_range6704w6706w & wire_y_pipeff_8_w_lg_w_q_range6704w6706w & wire_y_pipeff_8_w_lg_w_q_range6704w6706w & wire_y_pipeff_8_w_lg_w_q_range6704w6706w & wire_y_pipeff_8_w_lg_w_q_range6704w6706w & wire_y_pipeff_8_w_lg_w_q_range6704w6706w & wire_y_pipeff_8_w_lg_w_q_range6704w6706w & wire_y_pipeff_8_w_lg_w_q_range6890w6892w & wire_y_pipeff_8_w_lg_w_q_range6884w6886w & wire_y_pipeff_8_w_lg_w_q_range6878w6880w & wire_y_pipeff_8_w_lg_w_q_range6872w6874w & wire_y_pipeff_8_w_lg_w_q_range6866w6868w & wire_y_pipeff_8_w_lg_w_q_range6860w6862w & wire_y_pipeff_8_w_lg_w_q_range6854w6856w & wire_y_pipeff_8_w_lg_w_q_range6848w6850w & wire_y_pipeff_8_w_lg_w_q_range6842w6844w & wire_y_pipeff_8_w_lg_w_q_range6836w6838w & wire_y_pipeff_8_w_lg_w_q_range6830w6832w & wire_y_pipeff_8_w_lg_w_q_range6824w6826w & wire_y_pipeff_8_w_lg_w_q_range6818w6820w & wire_y_pipeff_8_w_lg_w_q_range6812w6814w & wire_y_pipeff_8_w_lg_w_q_range6806w6808w & wire_y_pipeff_8_w_lg_w_q_range6800w6802w & wire_y_pipeff_8_w_lg_w_q_range6794w6796w & wire_y_pipeff_8_w_lg_w_q_range6788w6790w & wire_y_pipeff_8_w_lg_w_q_range6782w6784w & wire_y_pipeff_8_w_lg_w_q_range6776w6778w & wire_y_pipeff_8_w_lg_w_q_range6770w6772w & wire_y_pipeff_8_w_lg_w_q_range6764w6766w & wire_y_pipeff_8_w_lg_w_q_range6758w6760w & wire_y_pipeff_8_w_lg_w_q_range6752w6754w & wire_y_pipeff_8_w_lg_w_q_range6747w6749w);
	x_prenodetwo_10_w <= ( wire_y_pipeff_9_w_lg_w_q_range7521w7523w & wire_y_pipeff_9_w_lg_w_q_range7521w7523w & wire_y_pipeff_9_w_lg_w_q_range7521w7523w & wire_y_pipeff_9_w_lg_w_q_range7521w7523w & wire_y_pipeff_9_w_lg_w_q_range7521w7523w & wire_y_pipeff_9_w_lg_w_q_range7521w7523w & wire_y_pipeff_9_w_lg_w_q_range7521w7523w & wire_y_pipeff_9_w_lg_w_q_range7521w7523w & wire_y_pipeff_9_w_lg_w_q_range7521w7523w & wire_y_pipeff_9_w_lg_w_q_range7521w7523w & wire_y_pipeff_9_w_lg_w_q_range7521w7523w & wire_y_pipeff_9_w_lg_w_q_range7521w7523w & wire_y_pipeff_9_w_lg_w_q_range7705w7707w & wire_y_pipeff_9_w_lg_w_q_range7699w7701w & wire_y_pipeff_9_w_lg_w_q_range7693w7695w & wire_y_pipeff_9_w_lg_w_q_range7687w7689w & wire_y_pipeff_9_w_lg_w_q_range7681w7683w & wire_y_pipeff_9_w_lg_w_q_range7675w7677w & wire_y_pipeff_9_w_lg_w_q_range7669w7671w & wire_y_pipeff_9_w_lg_w_q_range7663w7665w & wire_y_pipeff_9_w_lg_w_q_range7657w7659w & wire_y_pipeff_9_w_lg_w_q_range7651w7653w & wire_y_pipeff_9_w_lg_w_q_range7645w7647w & wire_y_pipeff_9_w_lg_w_q_range7639w7641w & wire_y_pipeff_9_w_lg_w_q_range7633w7635w & wire_y_pipeff_9_w_lg_w_q_range7627w7629w & wire_y_pipeff_9_w_lg_w_q_range7621w7623w & wire_y_pipeff_9_w_lg_w_q_range7615w7617w & wire_y_pipeff_9_w_lg_w_q_range7609w7611w & wire_y_pipeff_9_w_lg_w_q_range7603w7605w & wire_y_pipeff_9_w_lg_w_q_range7597w7599w & wire_y_pipeff_9_w_lg_w_q_range7591w7593w & wire_y_pipeff_9_w_lg_w_q_range7585w7587w & wire_y_pipeff_9_w_lg_w_q_range7579w7581w);
	x_prenodetwo_11_w <= ( wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8333w8335w & wire_y_pipeff_10_w_lg_w_q_range8515w8517w & wire_y_pipeff_10_w_lg_w_q_range8509w8511w & wire_y_pipeff_10_w_lg_w_q_range8503w8505w & wire_y_pipeff_10_w_lg_w_q_range8497w8499w & wire_y_pipeff_10_w_lg_w_q_range8491w8493w & wire_y_pipeff_10_w_lg_w_q_range8485w8487w & wire_y_pipeff_10_w_lg_w_q_range8479w8481w & wire_y_pipeff_10_w_lg_w_q_range8473w8475w & wire_y_pipeff_10_w_lg_w_q_range8467w8469w & wire_y_pipeff_10_w_lg_w_q_range8461w8463w & wire_y_pipeff_10_w_lg_w_q_range8455w8457w & wire_y_pipeff_10_w_lg_w_q_range8449w8451w & wire_y_pipeff_10_w_lg_w_q_range8443w8445w & wire_y_pipeff_10_w_lg_w_q_range8437w8439w & wire_y_pipeff_10_w_lg_w_q_range8431w8433w & wire_y_pipeff_10_w_lg_w_q_range8425w8427w & wire_y_pipeff_10_w_lg_w_q_range8419w8421w & wire_y_pipeff_10_w_lg_w_q_range8413w8415w & wire_y_pipeff_10_w_lg_w_q_range8407w8409w & wire_y_pipeff_10_w_lg_w_q_range8401w8403w & wire_y_pipeff_10_w_lg_w_q_range8395w8397w);
	x_prenodetwo_12_w <= ( wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9140w9142w & wire_y_pipeff_11_w_lg_w_q_range9320w9322w & wire_y_pipeff_11_w_lg_w_q_range9314w9316w & wire_y_pipeff_11_w_lg_w_q_range9308w9310w & wire_y_pipeff_11_w_lg_w_q_range9302w9304w & wire_y_pipeff_11_w_lg_w_q_range9296w9298w & wire_y_pipeff_11_w_lg_w_q_range9290w9292w & wire_y_pipeff_11_w_lg_w_q_range9284w9286w & wire_y_pipeff_11_w_lg_w_q_range9278w9280w & wire_y_pipeff_11_w_lg_w_q_range9272w9274w & wire_y_pipeff_11_w_lg_w_q_range9266w9268w & wire_y_pipeff_11_w_lg_w_q_range9260w9262w & wire_y_pipeff_11_w_lg_w_q_range9254w9256w & wire_y_pipeff_11_w_lg_w_q_range9248w9250w & wire_y_pipeff_11_w_lg_w_q_range9242w9244w & wire_y_pipeff_11_w_lg_w_q_range9236w9238w & wire_y_pipeff_11_w_lg_w_q_range9230w9232w & wire_y_pipeff_11_w_lg_w_q_range9224w9226w & wire_y_pipeff_11_w_lg_w_q_range9218w9220w & wire_y_pipeff_11_w_lg_w_q_range9212w9214w & wire_y_pipeff_11_w_lg_w_q_range9206w9208w);
	x_prenodetwo_13_w <= ( wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range9942w9944w & wire_y_pipeff_12_w_lg_w_q_range10120w10122w & wire_y_pipeff_12_w_lg_w_q_range10114w10116w & wire_y_pipeff_12_w_lg_w_q_range10108w10110w & wire_y_pipeff_12_w_lg_w_q_range10102w10104w & wire_y_pipeff_12_w_lg_w_q_range10096w10098w & wire_y_pipeff_12_w_lg_w_q_range10090w10092w & wire_y_pipeff_12_w_lg_w_q_range10084w10086w & wire_y_pipeff_12_w_lg_w_q_range10078w10080w & wire_y_pipeff_12_w_lg_w_q_range10072w10074w & wire_y_pipeff_12_w_lg_w_q_range10066w10068w & wire_y_pipeff_12_w_lg_w_q_range10060w10062w & wire_y_pipeff_12_w_lg_w_q_range10054w10056w & wire_y_pipeff_12_w_lg_w_q_range10048w10050w & wire_y_pipeff_12_w_lg_w_q_range10042w10044w & wire_y_pipeff_12_w_lg_w_q_range10036w10038w & wire_y_pipeff_12_w_lg_w_q_range10030w10032w & wire_y_pipeff_12_w_lg_w_q_range10024w10026w & wire_y_pipeff_12_w_lg_w_q_range10018w10020w & wire_y_pipeff_12_w_lg_w_q_range10012w10014w);
	x_prenodetwo_2_w <= ( wire_y_pipeff_1_w_lg_w_q_range845w847w & wire_y_pipeff_1_w_lg_w_q_range845w847w & wire_y_pipeff_1_w_lg_w_q_range845w847w & wire_y_pipeff_1_w_lg_w_q_range845w847w & wire_y_pipeff_1_w_lg_w_q_range1045w1047w & wire_y_pipeff_1_w_lg_w_q_range1039w1041w & wire_y_pipeff_1_w_lg_w_q_range1033w1035w & wire_y_pipeff_1_w_lg_w_q_range1027w1029w & wire_y_pipeff_1_w_lg_w_q_range1021w1023w & wire_y_pipeff_1_w_lg_w_q_range1015w1017w & wire_y_pipeff_1_w_lg_w_q_range1009w1011w & wire_y_pipeff_1_w_lg_w_q_range1003w1005w & wire_y_pipeff_1_w_lg_w_q_range997w999w & wire_y_pipeff_1_w_lg_w_q_range991w993w & wire_y_pipeff_1_w_lg_w_q_range985w987w & wire_y_pipeff_1_w_lg_w_q_range979w981w & wire_y_pipeff_1_w_lg_w_q_range973w975w & wire_y_pipeff_1_w_lg_w_q_range967w969w & wire_y_pipeff_1_w_lg_w_q_range961w963w & wire_y_pipeff_1_w_lg_w_q_range955w957w & wire_y_pipeff_1_w_lg_w_q_range949w951w & wire_y_pipeff_1_w_lg_w_q_range943w945w & wire_y_pipeff_1_w_lg_w_q_range937w939w & wire_y_pipeff_1_w_lg_w_q_range931w933w & wire_y_pipeff_1_w_lg_w_q_range925w927w & wire_y_pipeff_1_w_lg_w_q_range919w921w & wire_y_pipeff_1_w_lg_w_q_range913w915w & wire_y_pipeff_1_w_lg_w_q_range907w909w & wire_y_pipeff_1_w_lg_w_q_range901w903w & wire_y_pipeff_1_w_lg_w_q_range895w897w & wire_y_pipeff_1_w_lg_w_q_range889w891w & wire_y_pipeff_1_w_lg_w_q_range883w885w & wire_y_pipeff_1_w_lg_w_q_range877w879w & wire_y_pipeff_1_w_lg_w_q_range871w873w);
	x_prenodetwo_3_w <= ( wire_y_pipeff_2_w_lg_w_q_range1697w1699w & wire_y_pipeff_2_w_lg_w_q_range1697w1699w & wire_y_pipeff_2_w_lg_w_q_range1697w1699w & wire_y_pipeff_2_w_lg_w_q_range1697w1699w & wire_y_pipeff_2_w_lg_w_q_range1697w1699w & wire_y_pipeff_2_w_lg_w_q_range1895w1897w & wire_y_pipeff_2_w_lg_w_q_range1889w1891w & wire_y_pipeff_2_w_lg_w_q_range1883w1885w & wire_y_pipeff_2_w_lg_w_q_range1877w1879w & wire_y_pipeff_2_w_lg_w_q_range1871w1873w & wire_y_pipeff_2_w_lg_w_q_range1865w1867w & wire_y_pipeff_2_w_lg_w_q_range1859w1861w & wire_y_pipeff_2_w_lg_w_q_range1853w1855w & wire_y_pipeff_2_w_lg_w_q_range1847w1849w & wire_y_pipeff_2_w_lg_w_q_range1841w1843w & wire_y_pipeff_2_w_lg_w_q_range1835w1837w & wire_y_pipeff_2_w_lg_w_q_range1829w1831w & wire_y_pipeff_2_w_lg_w_q_range1823w1825w & wire_y_pipeff_2_w_lg_w_q_range1817w1819w & wire_y_pipeff_2_w_lg_w_q_range1811w1813w & wire_y_pipeff_2_w_lg_w_q_range1805w1807w & wire_y_pipeff_2_w_lg_w_q_range1799w1801w & wire_y_pipeff_2_w_lg_w_q_range1793w1795w & wire_y_pipeff_2_w_lg_w_q_range1787w1789w & wire_y_pipeff_2_w_lg_w_q_range1781w1783w & wire_y_pipeff_2_w_lg_w_q_range1775w1777w & wire_y_pipeff_2_w_lg_w_q_range1769w1771w & wire_y_pipeff_2_w_lg_w_q_range1763w1765w & wire_y_pipeff_2_w_lg_w_q_range1757w1759w & wire_y_pipeff_2_w_lg_w_q_range1751w1753w & wire_y_pipeff_2_w_lg_w_q_range1745w1747w & wire_y_pipeff_2_w_lg_w_q_range1739w1741w & wire_y_pipeff_2_w_lg_w_q_range1733w1735w & wire_y_pipeff_2_w_lg_w_q_range1727w1729w);
	x_prenodetwo_4_w <= ( wire_y_pipeff_3_w_lg_w_q_range2544w2546w & wire_y_pipeff_3_w_lg_w_q_range2544w2546w & wire_y_pipeff_3_w_lg_w_q_range2544w2546w & wire_y_pipeff_3_w_lg_w_q_range2544w2546w & wire_y_pipeff_3_w_lg_w_q_range2544w2546w & wire_y_pipeff_3_w_lg_w_q_range2544w2546w & wire_y_pipeff_3_w_lg_w_q_range2740w2742w & wire_y_pipeff_3_w_lg_w_q_range2734w2736w & wire_y_pipeff_3_w_lg_w_q_range2728w2730w & wire_y_pipeff_3_w_lg_w_q_range2722w2724w & wire_y_pipeff_3_w_lg_w_q_range2716w2718w & wire_y_pipeff_3_w_lg_w_q_range2710w2712w & wire_y_pipeff_3_w_lg_w_q_range2704w2706w & wire_y_pipeff_3_w_lg_w_q_range2698w2700w & wire_y_pipeff_3_w_lg_w_q_range2692w2694w & wire_y_pipeff_3_w_lg_w_q_range2686w2688w & wire_y_pipeff_3_w_lg_w_q_range2680w2682w & wire_y_pipeff_3_w_lg_w_q_range2674w2676w & wire_y_pipeff_3_w_lg_w_q_range2668w2670w & wire_y_pipeff_3_w_lg_w_q_range2662w2664w & wire_y_pipeff_3_w_lg_w_q_range2656w2658w & wire_y_pipeff_3_w_lg_w_q_range2650w2652w & wire_y_pipeff_3_w_lg_w_q_range2644w2646w & wire_y_pipeff_3_w_lg_w_q_range2638w2640w & wire_y_pipeff_3_w_lg_w_q_range2632w2634w & wire_y_pipeff_3_w_lg_w_q_range2626w2628w & wire_y_pipeff_3_w_lg_w_q_range2620w2622w & wire_y_pipeff_3_w_lg_w_q_range2614w2616w & wire_y_pipeff_3_w_lg_w_q_range2608w2610w & wire_y_pipeff_3_w_lg_w_q_range2602w2604w & wire_y_pipeff_3_w_lg_w_q_range2596w2598w & wire_y_pipeff_3_w_lg_w_q_range2590w2592w & wire_y_pipeff_3_w_lg_w_q_range2584w2586w & wire_y_pipeff_3_w_lg_w_q_range2578w2580w);
	x_prenodetwo_5_w <= ( wire_y_pipeff_4_w_lg_w_q_range3386w3388w & wire_y_pipeff_4_w_lg_w_q_range3386w3388w & wire_y_pipeff_4_w_lg_w_q_range3386w3388w & wire_y_pipeff_4_w_lg_w_q_range3386w3388w & wire_y_pipeff_4_w_lg_w_q_range3386w3388w & wire_y_pipeff_4_w_lg_w_q_range3386w3388w & wire_y_pipeff_4_w_lg_w_q_range3386w3388w & wire_y_pipeff_4_w_lg_w_q_range3580w3582w & wire_y_pipeff_4_w_lg_w_q_range3574w3576w & wire_y_pipeff_4_w_lg_w_q_range3568w3570w & wire_y_pipeff_4_w_lg_w_q_range3562w3564w & wire_y_pipeff_4_w_lg_w_q_range3556w3558w & wire_y_pipeff_4_w_lg_w_q_range3550w3552w & wire_y_pipeff_4_w_lg_w_q_range3544w3546w & wire_y_pipeff_4_w_lg_w_q_range3538w3540w & wire_y_pipeff_4_w_lg_w_q_range3532w3534w & wire_y_pipeff_4_w_lg_w_q_range3526w3528w & wire_y_pipeff_4_w_lg_w_q_range3520w3522w & wire_y_pipeff_4_w_lg_w_q_range3514w3516w & wire_y_pipeff_4_w_lg_w_q_range3508w3510w & wire_y_pipeff_4_w_lg_w_q_range3502w3504w & wire_y_pipeff_4_w_lg_w_q_range3496w3498w & wire_y_pipeff_4_w_lg_w_q_range3490w3492w & wire_y_pipeff_4_w_lg_w_q_range3484w3486w & wire_y_pipeff_4_w_lg_w_q_range3478w3480w & wire_y_pipeff_4_w_lg_w_q_range3472w3474w & wire_y_pipeff_4_w_lg_w_q_range3466w3468w & wire_y_pipeff_4_w_lg_w_q_range3460w3462w & wire_y_pipeff_4_w_lg_w_q_range3454w3456w & wire_y_pipeff_4_w_lg_w_q_range3448w3450w & wire_y_pipeff_4_w_lg_w_q_range3442w3444w & wire_y_pipeff_4_w_lg_w_q_range3436w3438w & wire_y_pipeff_4_w_lg_w_q_range3430w3432w & wire_y_pipeff_4_w_lg_w_q_range3424w3426w);
	x_prenodetwo_6_w <= ( wire_y_pipeff_5_w_lg_w_q_range4223w4225w & wire_y_pipeff_5_w_lg_w_q_range4223w4225w & wire_y_pipeff_5_w_lg_w_q_range4223w4225w & wire_y_pipeff_5_w_lg_w_q_range4223w4225w & wire_y_pipeff_5_w_lg_w_q_range4223w4225w & wire_y_pipeff_5_w_lg_w_q_range4223w4225w & wire_y_pipeff_5_w_lg_w_q_range4223w4225w & wire_y_pipeff_5_w_lg_w_q_range4223w4225w & wire_y_pipeff_5_w_lg_w_q_range4415w4417w & wire_y_pipeff_5_w_lg_w_q_range4409w4411w & wire_y_pipeff_5_w_lg_w_q_range4403w4405w & wire_y_pipeff_5_w_lg_w_q_range4397w4399w & wire_y_pipeff_5_w_lg_w_q_range4391w4393w & wire_y_pipeff_5_w_lg_w_q_range4385w4387w & wire_y_pipeff_5_w_lg_w_q_range4379w4381w & wire_y_pipeff_5_w_lg_w_q_range4373w4375w & wire_y_pipeff_5_w_lg_w_q_range4367w4369w & wire_y_pipeff_5_w_lg_w_q_range4361w4363w & wire_y_pipeff_5_w_lg_w_q_range4355w4357w & wire_y_pipeff_5_w_lg_w_q_range4349w4351w & wire_y_pipeff_5_w_lg_w_q_range4343w4345w & wire_y_pipeff_5_w_lg_w_q_range4337w4339w & wire_y_pipeff_5_w_lg_w_q_range4331w4333w & wire_y_pipeff_5_w_lg_w_q_range4325w4327w & wire_y_pipeff_5_w_lg_w_q_range4319w4321w & wire_y_pipeff_5_w_lg_w_q_range4313w4315w & wire_y_pipeff_5_w_lg_w_q_range4307w4309w & wire_y_pipeff_5_w_lg_w_q_range4301w4303w & wire_y_pipeff_5_w_lg_w_q_range4295w4297w & wire_y_pipeff_5_w_lg_w_q_range4289w4291w & wire_y_pipeff_5_w_lg_w_q_range4283w4285w & wire_y_pipeff_5_w_lg_w_q_range4277w4279w & wire_y_pipeff_5_w_lg_w_q_range4271w4273w & wire_y_pipeff_5_w_lg_w_q_range4265w4267w);
	x_prenodetwo_7_w <= ( wire_y_pipeff_6_w_lg_w_q_range5055w5057w & wire_y_pipeff_6_w_lg_w_q_range5055w5057w & wire_y_pipeff_6_w_lg_w_q_range5055w5057w & wire_y_pipeff_6_w_lg_w_q_range5055w5057w & wire_y_pipeff_6_w_lg_w_q_range5055w5057w & wire_y_pipeff_6_w_lg_w_q_range5055w5057w & wire_y_pipeff_6_w_lg_w_q_range5055w5057w & wire_y_pipeff_6_w_lg_w_q_range5055w5057w & wire_y_pipeff_6_w_lg_w_q_range5055w5057w & wire_y_pipeff_6_w_lg_w_q_range5245w5247w & wire_y_pipeff_6_w_lg_w_q_range5239w5241w & wire_y_pipeff_6_w_lg_w_q_range5233w5235w & wire_y_pipeff_6_w_lg_w_q_range5227w5229w & wire_y_pipeff_6_w_lg_w_q_range5221w5223w & wire_y_pipeff_6_w_lg_w_q_range5215w5217w & wire_y_pipeff_6_w_lg_w_q_range5209w5211w & wire_y_pipeff_6_w_lg_w_q_range5203w5205w & wire_y_pipeff_6_w_lg_w_q_range5197w5199w & wire_y_pipeff_6_w_lg_w_q_range5191w5193w & wire_y_pipeff_6_w_lg_w_q_range5185w5187w & wire_y_pipeff_6_w_lg_w_q_range5179w5181w & wire_y_pipeff_6_w_lg_w_q_range5173w5175w & wire_y_pipeff_6_w_lg_w_q_range5167w5169w & wire_y_pipeff_6_w_lg_w_q_range5161w5163w & wire_y_pipeff_6_w_lg_w_q_range5155w5157w & wire_y_pipeff_6_w_lg_w_q_range5149w5151w & wire_y_pipeff_6_w_lg_w_q_range5143w5145w & wire_y_pipeff_6_w_lg_w_q_range5137w5139w & wire_y_pipeff_6_w_lg_w_q_range5131w5133w & wire_y_pipeff_6_w_lg_w_q_range5125w5127w & wire_y_pipeff_6_w_lg_w_q_range5119w5121w & wire_y_pipeff_6_w_lg_w_q_range5113w5115w & wire_y_pipeff_6_w_lg_w_q_range5107w5109w & wire_y_pipeff_6_w_lg_w_q_range5101w5103w);
	x_prenodetwo_8_w <= ( wire_y_pipeff_7_w_lg_w_q_range5882w5884w & wire_y_pipeff_7_w_lg_w_q_range5882w5884w & wire_y_pipeff_7_w_lg_w_q_range5882w5884w & wire_y_pipeff_7_w_lg_w_q_range5882w5884w & wire_y_pipeff_7_w_lg_w_q_range5882w5884w & wire_y_pipeff_7_w_lg_w_q_range5882w5884w & wire_y_pipeff_7_w_lg_w_q_range5882w5884w & wire_y_pipeff_7_w_lg_w_q_range5882w5884w & wire_y_pipeff_7_w_lg_w_q_range5882w5884w & wire_y_pipeff_7_w_lg_w_q_range5882w5884w & wire_y_pipeff_7_w_lg_w_q_range6070w6072w & wire_y_pipeff_7_w_lg_w_q_range6064w6066w & wire_y_pipeff_7_w_lg_w_q_range6058w6060w & wire_y_pipeff_7_w_lg_w_q_range6052w6054w & wire_y_pipeff_7_w_lg_w_q_range6046w6048w & wire_y_pipeff_7_w_lg_w_q_range6040w6042w & wire_y_pipeff_7_w_lg_w_q_range6034w6036w & wire_y_pipeff_7_w_lg_w_q_range6028w6030w & wire_y_pipeff_7_w_lg_w_q_range6022w6024w & wire_y_pipeff_7_w_lg_w_q_range6016w6018w & wire_y_pipeff_7_w_lg_w_q_range6010w6012w & wire_y_pipeff_7_w_lg_w_q_range6004w6006w & wire_y_pipeff_7_w_lg_w_q_range5998w6000w & wire_y_pipeff_7_w_lg_w_q_range5992w5994w & wire_y_pipeff_7_w_lg_w_q_range5986w5988w & wire_y_pipeff_7_w_lg_w_q_range5980w5982w & wire_y_pipeff_7_w_lg_w_q_range5974w5976w & wire_y_pipeff_7_w_lg_w_q_range5968w5970w & wire_y_pipeff_7_w_lg_w_q_range5962w5964w & wire_y_pipeff_7_w_lg_w_q_range5956w5958w & wire_y_pipeff_7_w_lg_w_q_range5950w5952w & wire_y_pipeff_7_w_lg_w_q_range5944w5946w & wire_y_pipeff_7_w_lg_w_q_range5938w5940w & wire_y_pipeff_7_w_lg_w_q_range5932w5934w);
	x_prenodetwo_9_w <= ( wire_y_pipeff_8_w_lg_w_q_range6704w6706w & wire_y_pipeff_8_w_lg_w_q_range6704w6706w & wire_y_pipeff_8_w_lg_w_q_range6704w6706w & wire_y_pipeff_8_w_lg_w_q_range6704w6706w & wire_y_pipeff_8_w_lg_w_q_range6704w6706w & wire_y_pipeff_8_w_lg_w_q_range6704w6706w & wire_y_pipeff_8_w_lg_w_q_range6704w6706w & wire_y_pipeff_8_w_lg_w_q_range6704w6706w & wire_y_pipeff_8_w_lg_w_q_range6704w6706w & wire_y_pipeff_8_w_lg_w_q_range6704w6706w & wire_y_pipeff_8_w_lg_w_q_range6704w6706w & wire_y_pipeff_8_w_lg_w_q_range6890w6892w & wire_y_pipeff_8_w_lg_w_q_range6884w6886w & wire_y_pipeff_8_w_lg_w_q_range6878w6880w & wire_y_pipeff_8_w_lg_w_q_range6872w6874w & wire_y_pipeff_8_w_lg_w_q_range6866w6868w & wire_y_pipeff_8_w_lg_w_q_range6860w6862w & wire_y_pipeff_8_w_lg_w_q_range6854w6856w & wire_y_pipeff_8_w_lg_w_q_range6848w6850w & wire_y_pipeff_8_w_lg_w_q_range6842w6844w & wire_y_pipeff_8_w_lg_w_q_range6836w6838w & wire_y_pipeff_8_w_lg_w_q_range6830w6832w & wire_y_pipeff_8_w_lg_w_q_range6824w6826w & wire_y_pipeff_8_w_lg_w_q_range6818w6820w & wire_y_pipeff_8_w_lg_w_q_range6812w6814w & wire_y_pipeff_8_w_lg_w_q_range6806w6808w & wire_y_pipeff_8_w_lg_w_q_range6800w6802w & wire_y_pipeff_8_w_lg_w_q_range6794w6796w & wire_y_pipeff_8_w_lg_w_q_range6788w6790w & wire_y_pipeff_8_w_lg_w_q_range6782w6784w & wire_y_pipeff_8_w_lg_w_q_range6776w6778w & wire_y_pipeff_8_w_lg_w_q_range6770w6772w & wire_y_pipeff_8_w_lg_w_q_range6764w6766w & wire_y_pipeff_8_w_lg_w_q_range6758w6760w);
	x_start_node_w <= wire_cxs_value;
	x_subnode_10_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8049w8326w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8041w8318w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8033w8310w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8025w8302w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8017w8294w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8009w8286w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8001w8278w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7993w8270w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7985w8262w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7977w8254w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7969w8246w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7961w8238w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7953w8230w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7945w8222w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7937w8214w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7929w8206w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7921w8198w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7913w8190w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7905w8182w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7897w8174w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7889w8166w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7881w8158w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7873w8150w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7865w8142w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7857w8134w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7849w8126w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7841w8118w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7833w8110w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7825w8102w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7817w8094w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7809w8086w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7801w8078w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7793w8070w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7782w8059w);
	x_subnode_11_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8856w9133w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8848w9125w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8840w9117w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8832w9109w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8824w9101w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8816w9093w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8808w9085w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8800w9077w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8792w9069w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8784w9061w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8776w9053w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8768w9045w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8760w9037w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8752w9029w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8744w9021w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8736w9013w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8728w9005w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8720w8997w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8712w8989w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8704w8981w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8696w8973w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8688w8965w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8680w8957w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8672w8949w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8664w8941w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8656w8933w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8648w8925w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8640w8917w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8632w8909w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8624w8901w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8616w8893w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8608w8885w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8600w8877w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8589w8866w);
	x_subnode_12_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9658w9935w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9650w9927w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9642w9919w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9634w9911w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9626w9903w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9618w9895w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9610w9887w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9602w9879w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9594w9871w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9586w9863w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9578w9855w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9570w9847w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9562w9839w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9554w9831w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9546w9823w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9538w9815w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9530w9807w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9522w9799w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9514w9791w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9506w9783w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9498w9775w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9490w9767w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9482w9759w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9474w9751w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9466w9743w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9458w9735w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9450w9727w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9442w9719w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9434w9711w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9426w9703w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9418w9695w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9410w9687w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9402w9679w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9391w9668w);
	x_subnode_13_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10455w10732w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10447w10724w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10439w10716w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10431w10708w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10423w10700w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10415w10692w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10407w10684w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10399w10676w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10391w10668w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10383w10660w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10375w10652w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10367w10644w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10359w10636w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10351w10628w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10343w10620w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10335w10612w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10327w10604w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10319w10596w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10311w10588w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10303w10580w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10295w10572w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10287w10564w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10279w10556w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10271w10548w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10263w10540w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10255w10532w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10247w10524w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10239w10516w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10231w10508w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10223w10500w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10215w10492w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10207w10484w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10199w10476w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10188w10465w
);
	x_subnode_2_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1413w1690w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1405w1682w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1397w1674w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1389w1666w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1381w1658w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1373w1650w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1365w1642w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1357w1634w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1349w1626w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1341w1618w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1333w1610w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1325w1602w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1317w1594w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1309w1586w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1301w1578w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1293w1570w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1285w1562w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1277w1554w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1269w1546w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1261w1538w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1253w1530w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1245w1522w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1237w1514w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1229w1506w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1221w1498w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1213w1490w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1205w1482w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1197w1474w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1189w1466w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1181w1458w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1173w1450w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1165w1442w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1157w1434w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1146w1423w);
	x_subnode_3_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2260w2537w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2252w2529w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2244w2521w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2236w2513w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2228w2505w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2220w2497w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2212w2489w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2204w2481w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2196w2473w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2188w2465w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2180w2457w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2172w2449w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2164w2441w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2156w2433w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2148w2425w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2140w2417w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2132w2409w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2124w2401w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2116w2393w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2108w2385w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2100w2377w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2092w2369w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2084w2361w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2076w2353w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2068w2345w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2060w2337w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2052w2329w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2044w2321w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2036w2313w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2028w2305w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2020w2297w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2012w2289w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2004w2281w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1993w2270w);
	x_subnode_4_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3102w3379w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3094w3371w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3086w3363w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3078w3355w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3070w3347w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3062w3339w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3054w3331w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3046w3323w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3038w3315w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3030w3307w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3022w3299w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3014w3291w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3006w3283w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2998w3275w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2990w3267w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2982w3259w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2974w3251w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2966w3243w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2958w3235w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2950w3227w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2942w3219w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2934w3211w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2926w3203w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2918w3195w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2910w3187w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2902w3179w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2894w3171w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2886w3163w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2878w3155w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2870w3147w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2862w3139w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2854w3131w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2846w3123w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2835w3112w);
	x_subnode_5_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3939w4216w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3931w4208w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3923w4200w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3915w4192w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3907w4184w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3899w4176w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3891w4168w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3883w4160w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3875w4152w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3867w4144w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3859w4136w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3851w4128w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3843w4120w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3835w4112w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3827w4104w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3819w4096w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3811w4088w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3803w4080w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3795w4072w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3787w4064w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3779w4056w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3771w4048w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3763w4040w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3755w4032w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3747w4024w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3739w4016w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3731w4008w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3723w4000w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3715w3992w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3707w3984w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3699w3976w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3691w3968w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3683w3960w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3672w3949w);
	x_subnode_6_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4771w5048w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4763w5040w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4755w5032w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4747w5024w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4739w5016w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4731w5008w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4723w5000w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4715w4992w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4707w4984w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4699w4976w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4691w4968w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4683w4960w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4675w4952w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4667w4944w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4659w4936w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4651w4928w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4643w4920w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4635w4912w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4627w4904w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4619w4896w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4611w4888w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4603w4880w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4595w4872w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4587w4864w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4579w4856w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4571w4848w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4563w4840w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4555w4832w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4547w4824w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4539w4816w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4531w4808w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4523w4800w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4515w4792w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4504w4781w);
	x_subnode_7_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5598w5875w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5590w5867w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5582w5859w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5574w5851w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5566w5843w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5558w5835w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5550w5827w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5542w5819w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5534w5811w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5526w5803w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5518w5795w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5510w5787w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5502w5779w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5494w5771w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5486w5763w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5478w5755w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5470w5747w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5462w5739w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5454w5731w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5446w5723w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5438w5715w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5430w5707w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5422w5699w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5414w5691w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5406w5683w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5398w5675w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5390w5667w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5382w5659w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5374w5651w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5366w5643w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5358w5635w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5350w5627w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5342w5619w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5331w5608w);
	x_subnode_8_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6420w6697w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6412w6689w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6404w6681w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6396w6673w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6388w6665w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6380w6657w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6372w6649w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6364w6641w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6356w6633w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6348w6625w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6340w6617w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6332w6609w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6324w6601w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6316w6593w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6308w6585w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6300w6577w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6292w6569w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6284w6561w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6276w6553w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6268w6545w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6260w6537w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6252w6529w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6244w6521w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6236w6513w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6228w6505w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6220w6497w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6212w6489w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6204w6481w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6196w6473w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6188w6465w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6180w6457w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6172w6449w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6164w6441w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6153w6430w);
	x_subnode_9_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7237w7514w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7229w7506w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7221w7498w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7213w7490w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7205w7482w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7197w7474w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7189w7466w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7181w7458w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7173w7450w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7165w7442w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7157w7434w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7149w7426w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7141w7418w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7133w7410w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7125w7402w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7117w7394w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7109w7386w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7101w7378w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7093w7370w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7085w7362w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7077w7354w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7069w7346w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7061w7338w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7053w7330w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7045w7322w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7037w7314w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7029w7306w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7021w7298w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7013w7290w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7005w7282w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6997w7274w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6989w7266w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6981w7258w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6970w7247w);
	y_pipenode_10_w <= wire_y_pipenode_10_add_result;
	y_pipenode_11_w <= wire_y_pipenode_11_add_result;
	y_pipenode_12_w <= wire_y_pipenode_12_add_result;
	y_pipenode_13_w <= wire_y_pipenode_13_add_result;
	y_pipenode_2_w <= wire_y_pipenode_2_add_result;
	y_pipenode_3_w <= wire_y_pipenode_3_add_result;
	y_pipenode_4_w <= wire_y_pipenode_4_add_result;
	y_pipenode_5_w <= wire_y_pipenode_5_add_result;
	y_pipenode_6_w <= wire_y_pipenode_6_add_result;
	y_pipenode_7_w <= wire_y_pipenode_7_add_result;
	y_pipenode_8_w <= wire_y_pipenode_8_add_result;
	y_pipenode_9_w <= wire_y_pipenode_9_add_result;
	y_prenode_10_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7543w8055w8056w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7541w8047w8048w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7539w8039w8040w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7537w8031w8032w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7535w8023w8024w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7533w8015w8016w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7531w8007w8008w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7529w7999w8000w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7526w7991w7992w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7712w7983w7984w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7709w7975w7976w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7703w7967w7968w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7697w7959w7960w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7691w7951w7952w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7685w7943w7944w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7679w7935w7936w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7673w7927w7928w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7667w7919w7920w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7661w7911w7912w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7655w7903w7904w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7649w7895w7896w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7643w7887w7888w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7637w7879w7880w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7631w7871w7872w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7625w7863w7864w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7619w7855w7856w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7613w7847w7848w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7607w7839w7840w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7601w7831w7832w
 & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7595w7823w7824w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7589w7815w7816w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7583w7807w7808w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7577w7799w7800w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7572w7790w7791w);
	y_prenode_11_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8357w8862w8863w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8355w8854w8855w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8353w8846w8847w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8351w8838w8839w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8349w8830w8831w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8347w8822w8823w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8345w8814w8815w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8343w8806w8807w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8341w8798w8799w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8338w8790w8791w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8522w8782w8783w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8519w8774w8775w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8513w8766w8767w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8507w8758w8759w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8501w8750w8751w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8495w8742w8743w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8489w8734w8735w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8483w8726w8727w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8477w8718w8719w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8471w8710w8711w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8465w8702w8703w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8459w8694w8695w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8453w8686w8687w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8447w8678w8679w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8441w8670w8671w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8435w8662w8663w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8429w8654w8655w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8423w8646w8647w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8417w8638w8639w
 & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8411w8630w8631w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8405w8622w8623w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8399w8614w8615w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8393w8606w8607w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8388w8597w8598w);
	y_prenode_12_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9166w9664w9665w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9164w9656w9657w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9162w9648w9649w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9160w9640w9641w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9158w9632w9633w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9156w9624w9625w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9154w9616w9617w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9152w9608w9609w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9150w9600w9601w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9148w9592w9593w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9145w9584w9585w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9327w9576w9577w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9324w9568w9569w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9318w9560w9561w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9312w9552w9553w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9306w9544w9545w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9300w9536w9537w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9294w9528w9529w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9288w9520w9521w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9282w9512w9513w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9276w9504w9505w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9270w9496w9497w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9264w9488w9489w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9258w9480w9481w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9252w9472w9473w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9246w9464w9465w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9240w9456w9457w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9234w9448w9449w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9228w9440w9441w
 & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9222w9432w9433w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9216w9424w9425w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9210w9416w9417w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9204w9408w9409w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9199w9399w9400w);
	y_prenode_13_w <= ( wire_ccc_cordic_m_w10462w & wire_ccc_cordic_m_w10454w & wire_ccc_cordic_m_w10446w & wire_ccc_cordic_m_w10438w & wire_ccc_cordic_m_w10430w & wire_ccc_cordic_m_w10422w & wire_ccc_cordic_m_w10414w & wire_ccc_cordic_m_w10406w & wire_ccc_cordic_m_w10398w & wire_ccc_cordic_m_w10390w & wire_ccc_cordic_m_w10382w & wire_ccc_cordic_m_w10374w & wire_ccc_cordic_m_w10366w & wire_ccc_cordic_m_w10358w & wire_ccc_cordic_m_w10350w & wire_ccc_cordic_m_w10342w & wire_ccc_cordic_m_w10334w & wire_ccc_cordic_m_w10326w & wire_ccc_cordic_m_w10318w & wire_ccc_cordic_m_w10310w & wire_ccc_cordic_m_w10302w & wire_ccc_cordic_m_w10294w & wire_ccc_cordic_m_w10286w & wire_ccc_cordic_m_w10278w & wire_ccc_cordic_m_w10270w & wire_ccc_cordic_m_w10262w & wire_ccc_cordic_m_w10254w & wire_ccc_cordic_m_w10246w & wire_ccc_cordic_m_w10238w & wire_ccc_cordic_m_w10230w & wire_ccc_cordic_m_w10222w & wire_ccc_cordic_m_w10214w & wire_ccc_cordic_m_w10206w & wire_ccc_cordic_m_w10197w);
	y_prenode_2_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range850w1419w1420w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1052w1411w1412w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1049w1403w1404w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1043w1395w1396w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1037w1387w1388w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1031w1379w1380w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1025w1371w1372w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1019w1363w1364w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1013w1355w1356w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1007w1347w1348w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1001w1339w1340w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range995w1331w1332w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range989w1323w1324w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range983w1315w1316w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range977w1307w1308w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range971w1299w1300w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range965w1291w1292w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range959w1283w1284w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range953w1275w1276w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range947w1267w1268w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range941w1259w1260w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range935w1251w1252w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range929w1243w1244w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range923w1235w1236w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range917w1227w1228w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range911w1219w1220w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range905w1211w1212w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range899w1203w1204w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range893w1195w1196w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range887w1187w1188w
 & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range881w1179w1180w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range875w1171w1172w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range869w1163w1164w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range864w1154w1155w);
	y_prenode_3_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1705w2266w2267w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1702w2258w2259w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1902w2250w2251w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1899w2242w2243w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1893w2234w2235w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1887w2226w2227w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1881w2218w2219w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1875w2210w2211w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1869w2202w2203w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1863w2194w2195w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1857w2186w2187w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1851w2178w2179w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1845w2170w2171w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1839w2162w2163w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1833w2154w2155w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1827w2146w2147w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1821w2138w2139w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1815w2130w2131w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1809w2122w2123w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1803w2114w2115w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1797w2106w2107w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1791w2098w2099w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1785w2090w2091w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1779w2082w2083w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1773w2074w2075w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1767w2066w2067w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1761w2058w2059w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1755w2050w2051w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1749w2042w2043w 
& wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1743w2034w2035w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1737w2026w2027w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1731w2018w2019w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1725w2010w2011w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1720w2001w2002w);
	y_prenode_4_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2554w3108w3109w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2552w3100w3101w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2549w3092w3093w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2747w3084w3085w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2744w3076w3077w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2738w3068w3069w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2732w3060w3061w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2726w3052w3053w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2720w3044w3045w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2714w3036w3037w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2708w3028w3029w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2702w3020w3021w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2696w3012w3013w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2690w3004w3005w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2684w2996w2997w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2678w2988w2989w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2672w2980w2981w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2666w2972w2973w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2660w2964w2965w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2654w2956w2957w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2648w2948w2949w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2642w2940w2941w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2636w2932w2933w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2630w2924w2925w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2624w2916w2917w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2618w2908w2909w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2612w2900w2901w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2606w2892w2893w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2600w2884w2885w 
& wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2594w2876w2877w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2588w2868w2869w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2582w2860w2861w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2576w2852w2853w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2571w2843w2844w);
	y_prenode_5_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3398w3945w3946w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3396w3937w3938w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3394w3929w3930w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3391w3921w3922w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3587w3913w3914w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3584w3905w3906w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3578w3897w3898w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3572w3889w3890w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3566w3881w3882w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3560w3873w3874w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3554w3865w3866w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3548w3857w3858w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3542w3849w3850w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3536w3841w3842w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3530w3833w3834w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3524w3825w3826w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3518w3817w3818w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3512w3809w3810w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3506w3801w3802w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3500w3793w3794w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3494w3785w3786w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3488w3777w3778w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3482w3769w3770w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3476w3761w3762w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3470w3753w3754w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3464w3745w3746w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3458w3737w3738w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3452w3729w3730w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3446w3721w3722w 
& wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3440w3713w3714w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3434w3705w3706w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3428w3697w3698w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3422w3689w3690w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3417w3680w3681w);
	y_prenode_6_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4237w4777w4778w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4235w4769w4770w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4233w4761w4762w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4231w4753w4754w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4228w4745w4746w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4422w4737w4738w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4419w4729w4730w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4413w4721w4722w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4407w4713w4714w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4401w4705w4706w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4395w4697w4698w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4389w4689w4690w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4383w4681w4682w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4377w4673w4674w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4371w4665w4666w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4365w4657w4658w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4359w4649w4650w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4353w4641w4642w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4347w4633w4634w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4341w4625w4626w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4335w4617w4618w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4329w4609w4610w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4323w4601w4602w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4317w4593w4594w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4311w4585w4586w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4305w4577w4578w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4299w4569w4570w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4293w4561w4562w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4287w4553w4554w 
& wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4281w4545w4546w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4275w4537w4538w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4269w4529w4530w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4263w4521w4522w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4258w4512w4513w);
	y_prenode_7_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5071w5604w5605w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5069w5596w5597w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5067w5588w5589w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5065w5580w5581w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5063w5572w5573w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5060w5564w5565w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5252w5556w5557w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5249w5548w5549w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5243w5540w5541w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5237w5532w5533w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5231w5524w5525w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5225w5516w5517w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5219w5508w5509w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5213w5500w5501w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5207w5492w5493w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5201w5484w5485w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5195w5476w5477w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5189w5468w5469w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5183w5460w5461w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5177w5452w5453w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5171w5444w5445w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5165w5436w5437w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5159w5428w5429w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5153w5420w5421w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5147w5412w5413w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5141w5404w5405w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5135w5396w5397w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5129w5388w5389w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5123w5380w5381w 
& wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5117w5372w5373w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5111w5364w5365w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5105w5356w5357w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5099w5348w5349w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5094w5339w5340w);
	y_prenode_8_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5900w6426w6427w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5898w6418w6419w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5896w6410w6411w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5894w6402w6403w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5892w6394w6395w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5890w6386w6387w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5887w6378w6379w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6077w6370w6371w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6074w6362w6363w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6068w6354w6355w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6062w6346w6347w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6056w6338w6339w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6050w6330w6331w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6044w6322w6323w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6038w6314w6315w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6032w6306w6307w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6026w6298w6299w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6020w6290w6291w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6014w6282w6283w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6008w6274w6275w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6002w6266w6267w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5996w6258w6259w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5990w6250w6251w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5984w6242w6243w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5978w6234w6235w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5972w6226w6227w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5966w6218w6219w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5960w6210w6211w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5954w6202w6203w 
& wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5948w6194w6195w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5942w6186w6187w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5936w6178w6179w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5930w6170w6171w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5925w6161w6162w);
	y_prenode_9_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6724w7243w7244w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6722w7235w7236w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6720w7227w7228w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6718w7219w7220w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6716w7211w7212w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6714w7203w7204w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6712w7195w7196w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6709w7187w7188w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6897w7179w7180w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6894w7171w7172w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6888w7163w7164w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6882w7155w7156w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6876w7147w7148w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6870w7139w7140w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6864w7131w7132w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6858w7123w7124w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6852w7115w7116w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6846w7107w7108w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6840w7099w7100w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6834w7091w7092w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6828w7083w7084w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6822w7075w7076w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6816w7067w7068w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6810w7059w7060w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6804w7051w7052w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6798w7043w7044w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6792w7035w7036w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6786w7027w7028w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6780w7019w7020w 
& wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6774w7011w7012w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6768w7003w7004w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6762w6995w6996w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6756w6987w6988w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6751w6978w6979w);
	y_prenodeone_10_w <= ( x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33 DOWNTO 9));
	y_prenodeone_11_w <= ( x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33 DOWNTO 10));
	y_prenodeone_12_w <= ( x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33 DOWNTO 11));
	y_prenodeone_13_w <= ( x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33 DOWNTO 12));
	y_prenodeone_2_w <= ( x_pipeff_1(33) & x_pipeff_1(33 DOWNTO 1));
	y_prenodeone_3_w <= ( x_pipeff_2(33) & x_pipeff_2(33) & x_pipeff_2(33 DOWNTO 2));
	y_prenodeone_4_w <= ( x_pipeff_3(33) & x_pipeff_3(33) & x_pipeff_3(33) & x_pipeff_3(33 DOWNTO 3));
	y_prenodeone_5_w <= ( x_pipeff_4(33) & x_pipeff_4(33) & x_pipeff_4(33) & x_pipeff_4(33) & x_pipeff_4(33 DOWNTO 4));
	y_prenodeone_6_w <= ( x_pipeff_5(33) & x_pipeff_5(33) & x_pipeff_5(33) & x_pipeff_5(33) & x_pipeff_5(33) & x_pipeff_5(33 DOWNTO 5));
	y_prenodeone_7_w <= ( x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33 DOWNTO 6));
	y_prenodeone_8_w <= ( x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33 DOWNTO 7));
	y_prenodeone_9_w <= ( x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33 DOWNTO 8));
	y_prenodetwo_10_w <= ( x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33 DOWNTO 11));
	y_prenodetwo_11_w <= ( x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33 DOWNTO 12));
	y_prenodetwo_12_w <= ( x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33 DOWNTO 13));
	y_prenodetwo_13_w <= ( x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33 DOWNTO 14));
	y_prenodetwo_2_w <= ( x_pipeff_1(33) & x_pipeff_1(33) & x_pipeff_1(33) & x_pipeff_1(33 DOWNTO 3));
	y_prenodetwo_3_w <= ( x_pipeff_2(33) & x_pipeff_2(33) & x_pipeff_2(33) & x_pipeff_2(33) & x_pipeff_2(33 DOWNTO 4));
	y_prenodetwo_4_w <= ( x_pipeff_3(33) & x_pipeff_3(33) & x_pipeff_3(33) & x_pipeff_3(33) & x_pipeff_3(33) & x_pipeff_3(33 DOWNTO 5));
	y_prenodetwo_5_w <= ( x_pipeff_4(33) & x_pipeff_4(33) & x_pipeff_4(33) & x_pipeff_4(33) & x_pipeff_4(33) & x_pipeff_4(33) & x_pipeff_4(33 DOWNTO 6));
	y_prenodetwo_6_w <= ( x_pipeff_5(33) & x_pipeff_5(33) & x_pipeff_5(33) & x_pipeff_5(33) & x_pipeff_5(33) & x_pipeff_5(33) & x_pipeff_5(33) & x_pipeff_5(33 DOWNTO 7));
	y_prenodetwo_7_w <= ( x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33 DOWNTO 8));
	y_prenodetwo_8_w <= ( x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33 DOWNTO 9));
	y_prenodetwo_9_w <= ( x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33 DOWNTO 10));
	y_subnode_10_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8053w8328w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8045w8320w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8037w8312w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8029w8304w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8021w8296w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8013w8288w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8005w8280w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7997w8272w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7989w8264w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7981w8256w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7973w8248w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7965w8240w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7957w8232w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7949w8224w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7941w8216w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7933w8208w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7925w8200w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7917w8192w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7909w8184w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7901w8176w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7893w8168w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7885w8160w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7877w8152w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7869w8144w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7861w8136w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7853w8128w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7845w8120w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7837w8112w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7829w8104w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7821w8096w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7813w8088w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7805w8080w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7797w8072w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7788w8062w);
	y_subnode_11_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8860w9135w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8852w9127w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8844w9119w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8836w9111w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8828w9103w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8820w9095w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8812w9087w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8804w9079w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8796w9071w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8788w9063w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8780w9055w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8772w9047w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8764w9039w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8756w9031w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8748w9023w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8740w9015w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8732w9007w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8724w8999w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8716w8991w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8708w8983w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8700w8975w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8692w8967w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8684w8959w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8676w8951w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8668w8943w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8660w8935w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8652w8927w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8644w8919w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8636w8911w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8628w8903w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8620w8895w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8612w8887w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8604w8879w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8595w8869w);
	y_subnode_12_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9662w9937w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9654w9929w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9646w9921w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9638w9913w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9630w9905w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9622w9897w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9614w9889w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9606w9881w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9598w9873w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9590w9865w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9582w9857w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9574w9849w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9566w9841w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9558w9833w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9550w9825w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9542w9817w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9534w9809w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9526w9801w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9518w9793w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9510w9785w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9502w9777w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9494w9769w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9486w9761w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9478w9753w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9470w9745w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9462w9737w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9454w9729w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9446w9721w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9438w9713w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9430w9705w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9422w9697w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9414w9689w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9406w9681w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9397w9671w);
	y_subnode_13_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10459w10734w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10451w10726w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10443w10718w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10435w10710w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10427w10702w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10419w10694w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10411w10686w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10403w10678w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10395w10670w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10387w10662w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10379w10654w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10371w10646w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10363w10638w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10355w10630w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10347w10622w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10339w10614w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10331w10606w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10323w10598w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10315w10590w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10307w10582w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10299w10574w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10291w10566w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10283w10558w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10275w10550w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10267w10542w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10259w10534w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10251w10526w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10243w10518w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10235w10510w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10227w10502w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10219w10494w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10211w10486w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10203w10478w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10194w10468w
);
	y_subnode_1_w <= ( wire_x_pipeff_0_w_lg_w_q_range836w844w & wire_x_pipeff_0_w_lg_w_q_range831w842w & wire_x_pipeff_0_w_lg_w_lg_w_q_range826w839w840w & wire_x_pipeff_0_w_lg_w_lg_w_q_range821w834w835w & wire_x_pipeff_0_w_lg_w_lg_w_q_range816w829w830w & wire_x_pipeff_0_w_lg_w_lg_w_q_range811w824w825w & wire_x_pipeff_0_w_lg_w_lg_w_q_range806w819w820w & wire_x_pipeff_0_w_lg_w_lg_w_q_range801w814w815w & wire_x_pipeff_0_w_lg_w_lg_w_q_range796w809w810w & wire_x_pipeff_0_w_lg_w_lg_w_q_range791w804w805w & wire_x_pipeff_0_w_lg_w_lg_w_q_range786w799w800w & wire_x_pipeff_0_w_lg_w_lg_w_q_range781w794w795w & wire_x_pipeff_0_w_lg_w_lg_w_q_range776w789w790w & wire_x_pipeff_0_w_lg_w_lg_w_q_range771w784w785w & wire_x_pipeff_0_w_lg_w_lg_w_q_range766w779w780w & wire_x_pipeff_0_w_lg_w_lg_w_q_range761w774w775w & wire_x_pipeff_0_w_lg_w_lg_w_q_range756w769w770w & wire_x_pipeff_0_w_lg_w_lg_w_q_range751w764w765w & wire_x_pipeff_0_w_lg_w_lg_w_q_range746w759w760w & wire_x_pipeff_0_w_lg_w_lg_w_q_range741w754w755w & wire_x_pipeff_0_w_lg_w_lg_w_q_range736w749w750w & wire_x_pipeff_0_w_lg_w_lg_w_q_range731w744w745w & wire_x_pipeff_0_w_lg_w_lg_w_q_range726w739w740w & wire_x_pipeff_0_w_lg_w_lg_w_q_range721w734w735w & wire_x_pipeff_0_w_lg_w_lg_w_q_range716w729w730w & wire_x_pipeff_0_w_lg_w_lg_w_q_range711w724w725w & wire_x_pipeff_0_w_lg_w_lg_w_q_range706w719w720w & wire_x_pipeff_0_w_lg_w_lg_w_q_range701w714w715w & wire_x_pipeff_0_w_lg_w_lg_w_q_range696w709w710w & wire_x_pipeff_0_w_lg_w_lg_w_q_range691w704w705w & wire_x_pipeff_0_w_lg_w_lg_w_q_range685w699w700w & wire_x_pipeff_0_w_lg_w_lg_w_q_range677w694w695w & wire_x_pipeff_0_w_lg_w_lg_w_q_range686w689w690w & wire_x_pipeff_0_w_lg_w_lg_w_q_range678w682w683w);
	y_subnode_2_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1417w1692w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1409w1684w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1401w1676w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1393w1668w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1385w1660w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1377w1652w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1369w1644w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1361w1636w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1353w1628w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1345w1620w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1337w1612w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1329w1604w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1321w1596w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1313w1588w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1305w1580w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1297w1572w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1289w1564w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1281w1556w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1273w1548w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1265w1540w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1257w1532w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1249w1524w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1241w1516w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1233w1508w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1225w1500w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1217w1492w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1209w1484w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1201w1476w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1193w1468w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1185w1460w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1177w1452w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1169w1444w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1161w1436w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1152w1426w);
	y_subnode_3_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2264w2539w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2256w2531w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2248w2523w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2240w2515w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2232w2507w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2224w2499w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2216w2491w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2208w2483w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2200w2475w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2192w2467w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2184w2459w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2176w2451w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2168w2443w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2160w2435w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2152w2427w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2144w2419w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2136w2411w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2128w2403w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2120w2395w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2112w2387w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2104w2379w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2096w2371w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2088w2363w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2080w2355w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2072w2347w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2064w2339w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2056w2331w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2048w2323w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2040w2315w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2032w2307w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2024w2299w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2016w2291w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2008w2283w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1999w2273w);
	y_subnode_4_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3106w3381w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3098w3373w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3090w3365w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3082w3357w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3074w3349w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3066w3341w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3058w3333w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3050w3325w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3042w3317w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3034w3309w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3026w3301w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3018w3293w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3010w3285w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3002w3277w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2994w3269w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2986w3261w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2978w3253w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2970w3245w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2962w3237w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2954w3229w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2946w3221w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2938w3213w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2930w3205w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2922w3197w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2914w3189w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2906w3181w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2898w3173w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2890w3165w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2882w3157w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2874w3149w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2866w3141w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2858w3133w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2850w3125w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2841w3115w);
	y_subnode_5_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3943w4218w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3935w4210w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3927w4202w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3919w4194w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3911w4186w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3903w4178w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3895w4170w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3887w4162w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3879w4154w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3871w4146w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3863w4138w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3855w4130w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3847w4122w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3839w4114w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3831w4106w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3823w4098w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3815w4090w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3807w4082w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3799w4074w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3791w4066w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3783w4058w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3775w4050w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3767w4042w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3759w4034w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3751w4026w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3743w4018w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3735w4010w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3727w4002w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3719w3994w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3711w3986w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3703w3978w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3695w3970w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3687w3962w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3678w3952w);
	y_subnode_6_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4775w5050w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4767w5042w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4759w5034w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4751w5026w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4743w5018w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4735w5010w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4727w5002w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4719w4994w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4711w4986w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4703w4978w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4695w4970w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4687w4962w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4679w4954w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4671w4946w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4663w4938w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4655w4930w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4647w4922w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4639w4914w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4631w4906w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4623w4898w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4615w4890w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4607w4882w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4599w4874w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4591w4866w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4583w4858w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4575w4850w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4567w4842w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4559w4834w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4551w4826w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4543w4818w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4535w4810w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4527w4802w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4519w4794w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4510w4784w);
	y_subnode_7_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5602w5877w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5594w5869w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5586w5861w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5578w5853w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5570w5845w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5562w5837w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5554w5829w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5546w5821w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5538w5813w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5530w5805w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5522w5797w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5514w5789w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5506w5781w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5498w5773w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5490w5765w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5482w5757w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5474w5749w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5466w5741w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5458w5733w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5450w5725w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5442w5717w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5434w5709w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5426w5701w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5418w5693w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5410w5685w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5402w5677w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5394w5669w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5386w5661w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5378w5653w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5370w5645w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5362w5637w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5354w5629w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5346w5621w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5337w5611w);
	y_subnode_8_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6424w6699w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6416w6691w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6408w6683w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6400w6675w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6392w6667w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6384w6659w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6376w6651w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6368w6643w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6360w6635w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6352w6627w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6344w6619w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6336w6611w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6328w6603w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6320w6595w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6312w6587w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6304w6579w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6296w6571w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6288w6563w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6280w6555w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6272w6547w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6264w6539w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6256w6531w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6248w6523w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6240w6515w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6232w6507w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6224w6499w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6216w6491w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6208w6483w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6200w6475w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6192w6467w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6184w6459w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6176w6451w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6168w6443w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6159w6433w);
	y_subnode_9_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7241w7516w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7233w7508w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7225w7500w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7217w7492w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7209w7484w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7201w7476w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7193w7468w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7185w7460w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7177w7452w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7169w7444w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7161w7436w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7153w7428w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7145w7420w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7137w7412w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7129w7404w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7121w7396w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7113w7388w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7105w7380w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7097w7372w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7089w7364w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7081w7356w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7073w7348w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7065w7340w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7057w7332w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7049w7324w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7041w7316w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7033w7308w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7025w7300w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7017w7292w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7009w7284w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7001w7276w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6993w7268w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6985w7260w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6976w7250w);
	z_pipenode_10_w <= wire_z_pipenode_10_add_result;
	z_pipenode_11_w <= wire_z_pipenode_11_add_result;
	z_pipenode_12_w <= wire_z_pipenode_12_add_result;
	z_pipenode_13_w <= wire_z_pipenode_13_add_result;
	z_pipenode_2_w <= wire_z_pipenode_2_add_result;
	z_pipenode_3_w <= wire_z_pipenode_3_add_result;
	z_pipenode_4_w <= wire_z_pipenode_4_add_result;
	z_pipenode_5_w <= wire_z_pipenode_5_add_result;
	z_pipenode_6_w <= wire_z_pipenode_6_add_result;
	z_pipenode_7_w <= wire_z_pipenode_7_add_result;
	z_pipenode_8_w <= wire_z_pipenode_8_add_result;
	z_pipenode_9_w <= wire_z_pipenode_9_add_result;
	z_subnode_10_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8329w8331w8332w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8321w8323w8324w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8313w8315w8316w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8305w8307w8308w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8297w8299w8300w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8289w8291w8292w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8281w8283w8284w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8273w8275w8276w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8265w8267w8268w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8257w8259w8260w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8249w8251w8252w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8241w8243w8244w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8233w8235w8236w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8225w8227w8228w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8217w8219w8220w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8209w8211w8212w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8201w8203w8204w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8193w8195w8196w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8185w8187w8188w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8177w8179w8180w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8169w8171w8172w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8161w8163w8164w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8153w8155w8156w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8145w8147w8148w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8137w8139w8140w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8129w8131w8132w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8121w8123w8124w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8113w8115w8116w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8105w8107w8108w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8097w8099w8100w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8089w8091w8092w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8081w8083w8084w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8073w8075w8076w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8064w8066w8067w);
	z_subnode_11_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9136w9138w9139w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9128w9130w9131w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9120w9122w9123w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9112w9114w9115w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9104w9106w9107w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9096w9098w9099w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9088w9090w9091w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9080w9082w9083w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9072w9074w9075w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9064w9066w9067w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9056w9058w9059w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9048w9050w9051w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9040w9042w9043w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9032w9034w9035w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9024w9026w9027w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9016w9018w9019w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9008w9010w9011w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9000w9002w9003w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8992w8994w8995w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8984w8986w8987w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8976w8978w8979w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8968w8970w8971w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8960w8962w8963w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8952w8954w8955w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8944w8946w8947w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8936w8938w8939w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8928w8930w8931w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8920w8922w8923w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8912w8914w8915w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8904w8906w8907w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8896w8898w8899w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8888w8890w8891w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8880w8882w8883w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8871w8873w8874w);
	z_subnode_12_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9938w9940w9941w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9930w9932w9933w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9922w9924w9925w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9914w9916w9917w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9906w9908w9909w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9898w9900w9901w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9890w9892w9893w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9882w9884w9885w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9874w9876w9877w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9866w9868w9869w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9858w9860w9861w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9850w9852w9853w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9842w9844w9845w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9834w9836w9837w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9826w9828w9829w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9818w9820w9821w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9810w9812w9813w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9802w9804w9805w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9794w9796w9797w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9786w9788w9789w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9778w9780w9781w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9770w9772w9773w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9762w9764w9765w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9754w9756w9757w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9746w9748w9749w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9738w9740w9741w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9730w9732w9733w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9722w9724w9725w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9714w9716w9717w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9706w9708w9709w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9698w9700w9701w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9690w9692w9693w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9682w9684w9685w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9673w9675w9676w);
	z_subnode_13_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10735w10737w10738w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10727w10729w10730w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10719w10721w10722w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10711w10713w10714w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10703w10705w10706w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10695w10697w10698w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10687w10689w10690w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10679w10681w10682w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10671w10673w10674w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10663w10665w10666w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10655w10657w10658w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10647w10649w10650w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10639w10641w10642w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10631w10633w10634w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10623w10625w10626w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10615w10617w10618w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10607w10609w10610w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10599w10601w10602w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10591w10593w10594w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10583w10585w10586w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10575w10577w10578w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10567w10569w10570w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10559w10561w10562w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10551w10553w10554w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10543w10545w10546w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10535w10537w10538w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10527w10529w10530w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10519w10521w10522w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10511w10513w10514w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10503w10505w10506w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10495w10497w10498w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10487w10489w10490w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10479w10481w10482w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10470w10472w10473w);
	z_subnode_2_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1693w1695w1696w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1685w1687w1688w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1677w1679w1680w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1669w1671w1672w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1661w1663w1664w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1653w1655w1656w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1645w1647w1648w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1637w1639w1640w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1629w1631w1632w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1621w1623w1624w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1613w1615w1616w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1605w1607w1608w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1597w1599w1600w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1589w1591w1592w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1581w1583w1584w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1573w1575w1576w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1565w1567w1568w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1557w1559w1560w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1549w1551w1552w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1541w1543w1544w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1533w1535w1536w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1525w1527w1528w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1517w1519w1520w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1509w1511w1512w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1501w1503w1504w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1493w1495w1496w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1485w1487w1488w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1477w1479w1480w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1469w1471w1472w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1461w1463w1464w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1453w1455w1456w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1445w1447w1448w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1437w1439w1440w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1428w1430w1431w);
	z_subnode_3_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2540w2542w2543w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2532w2534w2535w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2524w2526w2527w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2516w2518w2519w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2508w2510w2511w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2500w2502w2503w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2492w2494w2495w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2484w2486w2487w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2476w2478w2479w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2468w2470w2471w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2460w2462w2463w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2452w2454w2455w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2444w2446w2447w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2436w2438w2439w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2428w2430w2431w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2420w2422w2423w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2412w2414w2415w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2404w2406w2407w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2396w2398w2399w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2388w2390w2391w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2380w2382w2383w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2372w2374w2375w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2364w2366w2367w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2356w2358w2359w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2348w2350w2351w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2340w2342w2343w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2332w2334w2335w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2324w2326w2327w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2316w2318w2319w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2308w2310w2311w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2300w2302w2303w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2292w2294w2295w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2284w2286w2287w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2275w2277w2278w);
	z_subnode_4_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3382w3384w3385w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3374w3376w3377w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3366w3368w3369w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3358w3360w3361w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3350w3352w3353w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3342w3344w3345w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3334w3336w3337w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3326w3328w3329w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3318w3320w3321w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3310w3312w3313w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3302w3304w3305w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3294w3296w3297w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3286w3288w3289w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3278w3280w3281w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3270w3272w3273w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3262w3264w3265w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3254w3256w3257w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3246w3248w3249w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3238w3240w3241w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3230w3232w3233w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3222w3224w3225w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3214w3216w3217w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3206w3208w3209w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3198w3200w3201w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3190w3192w3193w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3182w3184w3185w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3174w3176w3177w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3166w3168w3169w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3158w3160w3161w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3150w3152w3153w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3142w3144w3145w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3134w3136w3137w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3126w3128w3129w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3117w3119w3120w);
	z_subnode_5_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4219w4221w4222w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4211w4213w4214w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4203w4205w4206w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4195w4197w4198w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4187w4189w4190w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4179w4181w4182w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4171w4173w4174w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4163w4165w4166w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4155w4157w4158w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4147w4149w4150w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4139w4141w4142w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4131w4133w4134w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4123w4125w4126w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4115w4117w4118w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4107w4109w4110w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4099w4101w4102w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4091w4093w4094w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4083w4085w4086w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4075w4077w4078w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4067w4069w4070w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4059w4061w4062w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4051w4053w4054w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4043w4045w4046w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4035w4037w4038w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4027w4029w4030w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4019w4021w4022w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4011w4013w4014w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4003w4005w4006w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3995w3997w3998w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3987w3989w3990w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3979w3981w3982w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3971w3973w3974w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3963w3965w3966w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3954w3956w3957w);
	z_subnode_6_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5051w5053w5054w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5043w5045w5046w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5035w5037w5038w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5027w5029w5030w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5019w5021w5022w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5011w5013w5014w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5003w5005w5006w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4995w4997w4998w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4987w4989w4990w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4979w4981w4982w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4971w4973w4974w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4963w4965w4966w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4955w4957w4958w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4947w4949w4950w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4939w4941w4942w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4931w4933w4934w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4923w4925w4926w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4915w4917w4918w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4907w4909w4910w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4899w4901w4902w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4891w4893w4894w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4883w4885w4886w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4875w4877w4878w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4867w4869w4870w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4859w4861w4862w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4851w4853w4854w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4843w4845w4846w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4835w4837w4838w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4827w4829w4830w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4819w4821w4822w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4811w4813w4814w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4803w4805w4806w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4795w4797w4798w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4786w4788w4789w);
	z_subnode_7_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5878w5880w5881w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5870w5872w5873w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5862w5864w5865w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5854w5856w5857w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5846w5848w5849w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5838w5840w5841w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5830w5832w5833w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5822w5824w5825w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5814w5816w5817w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5806w5808w5809w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5798w5800w5801w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5790w5792w5793w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5782w5784w5785w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5774w5776w5777w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5766w5768w5769w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5758w5760w5761w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5750w5752w5753w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5742w5744w5745w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5734w5736w5737w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5726w5728w5729w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5718w5720w5721w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5710w5712w5713w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5702w5704w5705w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5694w5696w5697w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5686w5688w5689w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5678w5680w5681w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5670w5672w5673w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5662w5664w5665w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5654w5656w5657w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5646w5648w5649w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5638w5640w5641w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5630w5632w5633w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5622w5624w5625w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5613w5615w5616w);
	z_subnode_8_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6700w6702w6703w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6692w6694w6695w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6684w6686w6687w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6676w6678w6679w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6668w6670w6671w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6660w6662w6663w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6652w6654w6655w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6644w6646w6647w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6636w6638w6639w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6628w6630w6631w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6620w6622w6623w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6612w6614w6615w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6604w6606w6607w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6596w6598w6599w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6588w6590w6591w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6580w6582w6583w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6572w6574w6575w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6564w6566w6567w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6556w6558w6559w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6548w6550w6551w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6540w6542w6543w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6532w6534w6535w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6524w6526w6527w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6516w6518w6519w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6508w6510w6511w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6500w6502w6503w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6492w6494w6495w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6484w6486w6487w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6476w6478w6479w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6468w6470w6471w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6460w6462w6463w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6452w6454w6455w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6444w6446w6447w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6435w6437w6438w);
	z_subnode_9_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7517w7519w7520w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7509w7511w7512w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7501w7503w7504w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7493w7495w7496w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7485w7487w7488w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7477w7479w7480w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7469w7471w7472w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7461w7463w7464w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7453w7455w7456w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7445w7447w7448w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7437w7439w7440w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7429w7431w7432w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7421w7423w7424w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7413w7415w7416w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7405w7407w7408w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7397w7399w7400w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7389w7391w7392w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7381w7383w7384w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7373w7375w7376w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7365w7367w7368w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7357w7359w7360w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7349w7351w7352w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7341w7343w7344w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7333w7335w7336w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7325w7327w7328w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7317w7319w7320w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7309w7311w7312w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7301w7303w7304w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7293w7295w7296w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7285w7287w7288w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7277w7279w7280w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7269w7271w7272w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7261w7263w7264w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7252w7254w7255w);
	wire_ccc_cordic_m_w_atannode_10_w_range8871w(0) <= atannode_10_w(0);
	wire_ccc_cordic_m_w_atannode_10_w_range8952w(0) <= atannode_10_w(10);
	wire_ccc_cordic_m_w_atannode_10_w_range8960w(0) <= atannode_10_w(11);
	wire_ccc_cordic_m_w_atannode_10_w_range8968w(0) <= atannode_10_w(12);
	wire_ccc_cordic_m_w_atannode_10_w_range8976w(0) <= atannode_10_w(13);
	wire_ccc_cordic_m_w_atannode_10_w_range8984w(0) <= atannode_10_w(14);
	wire_ccc_cordic_m_w_atannode_10_w_range8992w(0) <= atannode_10_w(15);
	wire_ccc_cordic_m_w_atannode_10_w_range9000w(0) <= atannode_10_w(16);
	wire_ccc_cordic_m_w_atannode_10_w_range9008w(0) <= atannode_10_w(17);
	wire_ccc_cordic_m_w_atannode_10_w_range9016w(0) <= atannode_10_w(18);
	wire_ccc_cordic_m_w_atannode_10_w_range9024w(0) <= atannode_10_w(19);
	wire_ccc_cordic_m_w_atannode_10_w_range8880w(0) <= atannode_10_w(1);
	wire_ccc_cordic_m_w_atannode_10_w_range9032w(0) <= atannode_10_w(20);
	wire_ccc_cordic_m_w_atannode_10_w_range9040w(0) <= atannode_10_w(21);
	wire_ccc_cordic_m_w_atannode_10_w_range9048w(0) <= atannode_10_w(22);
	wire_ccc_cordic_m_w_atannode_10_w_range9056w(0) <= atannode_10_w(23);
	wire_ccc_cordic_m_w_atannode_10_w_range9064w(0) <= atannode_10_w(24);
	wire_ccc_cordic_m_w_atannode_10_w_range9072w(0) <= atannode_10_w(25);
	wire_ccc_cordic_m_w_atannode_10_w_range9080w(0) <= atannode_10_w(26);
	wire_ccc_cordic_m_w_atannode_10_w_range9088w(0) <= atannode_10_w(27);
	wire_ccc_cordic_m_w_atannode_10_w_range9096w(0) <= atannode_10_w(28);
	wire_ccc_cordic_m_w_atannode_10_w_range9104w(0) <= atannode_10_w(29);
	wire_ccc_cordic_m_w_atannode_10_w_range8888w(0) <= atannode_10_w(2);
	wire_ccc_cordic_m_w_atannode_10_w_range9112w(0) <= atannode_10_w(30);
	wire_ccc_cordic_m_w_atannode_10_w_range9120w(0) <= atannode_10_w(31);
	wire_ccc_cordic_m_w_atannode_10_w_range9128w(0) <= atannode_10_w(32);
	wire_ccc_cordic_m_w_atannode_10_w_range9136w(0) <= atannode_10_w(33);
	wire_ccc_cordic_m_w_atannode_10_w_range8896w(0) <= atannode_10_w(3);
	wire_ccc_cordic_m_w_atannode_10_w_range8904w(0) <= atannode_10_w(4);
	wire_ccc_cordic_m_w_atannode_10_w_range8912w(0) <= atannode_10_w(5);
	wire_ccc_cordic_m_w_atannode_10_w_range8920w(0) <= atannode_10_w(6);
	wire_ccc_cordic_m_w_atannode_10_w_range8928w(0) <= atannode_10_w(7);
	wire_ccc_cordic_m_w_atannode_10_w_range8936w(0) <= atannode_10_w(8);
	wire_ccc_cordic_m_w_atannode_10_w_range8944w(0) <= atannode_10_w(9);
	wire_ccc_cordic_m_w_atannode_11_w_range9673w(0) <= atannode_11_w(0);
	wire_ccc_cordic_m_w_atannode_11_w_range9754w(0) <= atannode_11_w(10);
	wire_ccc_cordic_m_w_atannode_11_w_range9762w(0) <= atannode_11_w(11);
	wire_ccc_cordic_m_w_atannode_11_w_range9770w(0) <= atannode_11_w(12);
	wire_ccc_cordic_m_w_atannode_11_w_range9778w(0) <= atannode_11_w(13);
	wire_ccc_cordic_m_w_atannode_11_w_range9786w(0) <= atannode_11_w(14);
	wire_ccc_cordic_m_w_atannode_11_w_range9794w(0) <= atannode_11_w(15);
	wire_ccc_cordic_m_w_atannode_11_w_range9802w(0) <= atannode_11_w(16);
	wire_ccc_cordic_m_w_atannode_11_w_range9810w(0) <= atannode_11_w(17);
	wire_ccc_cordic_m_w_atannode_11_w_range9818w(0) <= atannode_11_w(18);
	wire_ccc_cordic_m_w_atannode_11_w_range9826w(0) <= atannode_11_w(19);
	wire_ccc_cordic_m_w_atannode_11_w_range9682w(0) <= atannode_11_w(1);
	wire_ccc_cordic_m_w_atannode_11_w_range9834w(0) <= atannode_11_w(20);
	wire_ccc_cordic_m_w_atannode_11_w_range9842w(0) <= atannode_11_w(21);
	wire_ccc_cordic_m_w_atannode_11_w_range9850w(0) <= atannode_11_w(22);
	wire_ccc_cordic_m_w_atannode_11_w_range9858w(0) <= atannode_11_w(23);
	wire_ccc_cordic_m_w_atannode_11_w_range9866w(0) <= atannode_11_w(24);
	wire_ccc_cordic_m_w_atannode_11_w_range9874w(0) <= atannode_11_w(25);
	wire_ccc_cordic_m_w_atannode_11_w_range9882w(0) <= atannode_11_w(26);
	wire_ccc_cordic_m_w_atannode_11_w_range9890w(0) <= atannode_11_w(27);
	wire_ccc_cordic_m_w_atannode_11_w_range9898w(0) <= atannode_11_w(28);
	wire_ccc_cordic_m_w_atannode_11_w_range9906w(0) <= atannode_11_w(29);
	wire_ccc_cordic_m_w_atannode_11_w_range9690w(0) <= atannode_11_w(2);
	wire_ccc_cordic_m_w_atannode_11_w_range9914w(0) <= atannode_11_w(30);
	wire_ccc_cordic_m_w_atannode_11_w_range9922w(0) <= atannode_11_w(31);
	wire_ccc_cordic_m_w_atannode_11_w_range9930w(0) <= atannode_11_w(32);
	wire_ccc_cordic_m_w_atannode_11_w_range9938w(0) <= atannode_11_w(33);
	wire_ccc_cordic_m_w_atannode_11_w_range9698w(0) <= atannode_11_w(3);
	wire_ccc_cordic_m_w_atannode_11_w_range9706w(0) <= atannode_11_w(4);
	wire_ccc_cordic_m_w_atannode_11_w_range9714w(0) <= atannode_11_w(5);
	wire_ccc_cordic_m_w_atannode_11_w_range9722w(0) <= atannode_11_w(6);
	wire_ccc_cordic_m_w_atannode_11_w_range9730w(0) <= atannode_11_w(7);
	wire_ccc_cordic_m_w_atannode_11_w_range9738w(0) <= atannode_11_w(8);
	wire_ccc_cordic_m_w_atannode_11_w_range9746w(0) <= atannode_11_w(9);
	wire_ccc_cordic_m_w_atannode_12_w_range10470w(0) <= atannode_12_w(0);
	wire_ccc_cordic_m_w_atannode_12_w_range10551w(0) <= atannode_12_w(10);
	wire_ccc_cordic_m_w_atannode_12_w_range10559w(0) <= atannode_12_w(11);
	wire_ccc_cordic_m_w_atannode_12_w_range10567w(0) <= atannode_12_w(12);
	wire_ccc_cordic_m_w_atannode_12_w_range10575w(0) <= atannode_12_w(13);
	wire_ccc_cordic_m_w_atannode_12_w_range10583w(0) <= atannode_12_w(14);
	wire_ccc_cordic_m_w_atannode_12_w_range10591w(0) <= atannode_12_w(15);
	wire_ccc_cordic_m_w_atannode_12_w_range10599w(0) <= atannode_12_w(16);
	wire_ccc_cordic_m_w_atannode_12_w_range10607w(0) <= atannode_12_w(17);
	wire_ccc_cordic_m_w_atannode_12_w_range10615w(0) <= atannode_12_w(18);
	wire_ccc_cordic_m_w_atannode_12_w_range10623w(0) <= atannode_12_w(19);
	wire_ccc_cordic_m_w_atannode_12_w_range10479w(0) <= atannode_12_w(1);
	wire_ccc_cordic_m_w_atannode_12_w_range10631w(0) <= atannode_12_w(20);
	wire_ccc_cordic_m_w_atannode_12_w_range10639w(0) <= atannode_12_w(21);
	wire_ccc_cordic_m_w_atannode_12_w_range10647w(0) <= atannode_12_w(22);
	wire_ccc_cordic_m_w_atannode_12_w_range10655w(0) <= atannode_12_w(23);
	wire_ccc_cordic_m_w_atannode_12_w_range10663w(0) <= atannode_12_w(24);
	wire_ccc_cordic_m_w_atannode_12_w_range10671w(0) <= atannode_12_w(25);
	wire_ccc_cordic_m_w_atannode_12_w_range10679w(0) <= atannode_12_w(26);
	wire_ccc_cordic_m_w_atannode_12_w_range10687w(0) <= atannode_12_w(27);
	wire_ccc_cordic_m_w_atannode_12_w_range10695w(0) <= atannode_12_w(28);
	wire_ccc_cordic_m_w_atannode_12_w_range10703w(0) <= atannode_12_w(29);
	wire_ccc_cordic_m_w_atannode_12_w_range10487w(0) <= atannode_12_w(2);
	wire_ccc_cordic_m_w_atannode_12_w_range10711w(0) <= atannode_12_w(30);
	wire_ccc_cordic_m_w_atannode_12_w_range10719w(0) <= atannode_12_w(31);
	wire_ccc_cordic_m_w_atannode_12_w_range10727w(0) <= atannode_12_w(32);
	wire_ccc_cordic_m_w_atannode_12_w_range10735w(0) <= atannode_12_w(33);
	wire_ccc_cordic_m_w_atannode_12_w_range10495w(0) <= atannode_12_w(3);
	wire_ccc_cordic_m_w_atannode_12_w_range10503w(0) <= atannode_12_w(4);
	wire_ccc_cordic_m_w_atannode_12_w_range10511w(0) <= atannode_12_w(5);
	wire_ccc_cordic_m_w_atannode_12_w_range10519w(0) <= atannode_12_w(6);
	wire_ccc_cordic_m_w_atannode_12_w_range10527w(0) <= atannode_12_w(7);
	wire_ccc_cordic_m_w_atannode_12_w_range10535w(0) <= atannode_12_w(8);
	wire_ccc_cordic_m_w_atannode_12_w_range10543w(0) <= atannode_12_w(9);
	wire_ccc_cordic_m_w_atannode_1_w_range1428w(0) <= atannode_1_w(0);
	wire_ccc_cordic_m_w_atannode_1_w_range1509w(0) <= atannode_1_w(10);
	wire_ccc_cordic_m_w_atannode_1_w_range1517w(0) <= atannode_1_w(11);
	wire_ccc_cordic_m_w_atannode_1_w_range1525w(0) <= atannode_1_w(12);
	wire_ccc_cordic_m_w_atannode_1_w_range1533w(0) <= atannode_1_w(13);
	wire_ccc_cordic_m_w_atannode_1_w_range1541w(0) <= atannode_1_w(14);
	wire_ccc_cordic_m_w_atannode_1_w_range1549w(0) <= atannode_1_w(15);
	wire_ccc_cordic_m_w_atannode_1_w_range1557w(0) <= atannode_1_w(16);
	wire_ccc_cordic_m_w_atannode_1_w_range1565w(0) <= atannode_1_w(17);
	wire_ccc_cordic_m_w_atannode_1_w_range1573w(0) <= atannode_1_w(18);
	wire_ccc_cordic_m_w_atannode_1_w_range1581w(0) <= atannode_1_w(19);
	wire_ccc_cordic_m_w_atannode_1_w_range1437w(0) <= atannode_1_w(1);
	wire_ccc_cordic_m_w_atannode_1_w_range1589w(0) <= atannode_1_w(20);
	wire_ccc_cordic_m_w_atannode_1_w_range1597w(0) <= atannode_1_w(21);
	wire_ccc_cordic_m_w_atannode_1_w_range1605w(0) <= atannode_1_w(22);
	wire_ccc_cordic_m_w_atannode_1_w_range1613w(0) <= atannode_1_w(23);
	wire_ccc_cordic_m_w_atannode_1_w_range1621w(0) <= atannode_1_w(24);
	wire_ccc_cordic_m_w_atannode_1_w_range1629w(0) <= atannode_1_w(25);
	wire_ccc_cordic_m_w_atannode_1_w_range1637w(0) <= atannode_1_w(26);
	wire_ccc_cordic_m_w_atannode_1_w_range1645w(0) <= atannode_1_w(27);
	wire_ccc_cordic_m_w_atannode_1_w_range1653w(0) <= atannode_1_w(28);
	wire_ccc_cordic_m_w_atannode_1_w_range1661w(0) <= atannode_1_w(29);
	wire_ccc_cordic_m_w_atannode_1_w_range1445w(0) <= atannode_1_w(2);
	wire_ccc_cordic_m_w_atannode_1_w_range1669w(0) <= atannode_1_w(30);
	wire_ccc_cordic_m_w_atannode_1_w_range1677w(0) <= atannode_1_w(31);
	wire_ccc_cordic_m_w_atannode_1_w_range1685w(0) <= atannode_1_w(32);
	wire_ccc_cordic_m_w_atannode_1_w_range1693w(0) <= atannode_1_w(33);
	wire_ccc_cordic_m_w_atannode_1_w_range1453w(0) <= atannode_1_w(3);
	wire_ccc_cordic_m_w_atannode_1_w_range1461w(0) <= atannode_1_w(4);
	wire_ccc_cordic_m_w_atannode_1_w_range1469w(0) <= atannode_1_w(5);
	wire_ccc_cordic_m_w_atannode_1_w_range1477w(0) <= atannode_1_w(6);
	wire_ccc_cordic_m_w_atannode_1_w_range1485w(0) <= atannode_1_w(7);
	wire_ccc_cordic_m_w_atannode_1_w_range1493w(0) <= atannode_1_w(8);
	wire_ccc_cordic_m_w_atannode_1_w_range1501w(0) <= atannode_1_w(9);
	wire_ccc_cordic_m_w_atannode_2_w_range2275w(0) <= atannode_2_w(0);
	wire_ccc_cordic_m_w_atannode_2_w_range2356w(0) <= atannode_2_w(10);
	wire_ccc_cordic_m_w_atannode_2_w_range2364w(0) <= atannode_2_w(11);
	wire_ccc_cordic_m_w_atannode_2_w_range2372w(0) <= atannode_2_w(12);
	wire_ccc_cordic_m_w_atannode_2_w_range2380w(0) <= atannode_2_w(13);
	wire_ccc_cordic_m_w_atannode_2_w_range2388w(0) <= atannode_2_w(14);
	wire_ccc_cordic_m_w_atannode_2_w_range2396w(0) <= atannode_2_w(15);
	wire_ccc_cordic_m_w_atannode_2_w_range2404w(0) <= atannode_2_w(16);
	wire_ccc_cordic_m_w_atannode_2_w_range2412w(0) <= atannode_2_w(17);
	wire_ccc_cordic_m_w_atannode_2_w_range2420w(0) <= atannode_2_w(18);
	wire_ccc_cordic_m_w_atannode_2_w_range2428w(0) <= atannode_2_w(19);
	wire_ccc_cordic_m_w_atannode_2_w_range2284w(0) <= atannode_2_w(1);
	wire_ccc_cordic_m_w_atannode_2_w_range2436w(0) <= atannode_2_w(20);
	wire_ccc_cordic_m_w_atannode_2_w_range2444w(0) <= atannode_2_w(21);
	wire_ccc_cordic_m_w_atannode_2_w_range2452w(0) <= atannode_2_w(22);
	wire_ccc_cordic_m_w_atannode_2_w_range2460w(0) <= atannode_2_w(23);
	wire_ccc_cordic_m_w_atannode_2_w_range2468w(0) <= atannode_2_w(24);
	wire_ccc_cordic_m_w_atannode_2_w_range2476w(0) <= atannode_2_w(25);
	wire_ccc_cordic_m_w_atannode_2_w_range2484w(0) <= atannode_2_w(26);
	wire_ccc_cordic_m_w_atannode_2_w_range2492w(0) <= atannode_2_w(27);
	wire_ccc_cordic_m_w_atannode_2_w_range2500w(0) <= atannode_2_w(28);
	wire_ccc_cordic_m_w_atannode_2_w_range2508w(0) <= atannode_2_w(29);
	wire_ccc_cordic_m_w_atannode_2_w_range2292w(0) <= atannode_2_w(2);
	wire_ccc_cordic_m_w_atannode_2_w_range2516w(0) <= atannode_2_w(30);
	wire_ccc_cordic_m_w_atannode_2_w_range2524w(0) <= atannode_2_w(31);
	wire_ccc_cordic_m_w_atannode_2_w_range2532w(0) <= atannode_2_w(32);
	wire_ccc_cordic_m_w_atannode_2_w_range2540w(0) <= atannode_2_w(33);
	wire_ccc_cordic_m_w_atannode_2_w_range2300w(0) <= atannode_2_w(3);
	wire_ccc_cordic_m_w_atannode_2_w_range2308w(0) <= atannode_2_w(4);
	wire_ccc_cordic_m_w_atannode_2_w_range2316w(0) <= atannode_2_w(5);
	wire_ccc_cordic_m_w_atannode_2_w_range2324w(0) <= atannode_2_w(6);
	wire_ccc_cordic_m_w_atannode_2_w_range2332w(0) <= atannode_2_w(7);
	wire_ccc_cordic_m_w_atannode_2_w_range2340w(0) <= atannode_2_w(8);
	wire_ccc_cordic_m_w_atannode_2_w_range2348w(0) <= atannode_2_w(9);
	wire_ccc_cordic_m_w_atannode_3_w_range3117w(0) <= atannode_3_w(0);
	wire_ccc_cordic_m_w_atannode_3_w_range3198w(0) <= atannode_3_w(10);
	wire_ccc_cordic_m_w_atannode_3_w_range3206w(0) <= atannode_3_w(11);
	wire_ccc_cordic_m_w_atannode_3_w_range3214w(0) <= atannode_3_w(12);
	wire_ccc_cordic_m_w_atannode_3_w_range3222w(0) <= atannode_3_w(13);
	wire_ccc_cordic_m_w_atannode_3_w_range3230w(0) <= atannode_3_w(14);
	wire_ccc_cordic_m_w_atannode_3_w_range3238w(0) <= atannode_3_w(15);
	wire_ccc_cordic_m_w_atannode_3_w_range3246w(0) <= atannode_3_w(16);
	wire_ccc_cordic_m_w_atannode_3_w_range3254w(0) <= atannode_3_w(17);
	wire_ccc_cordic_m_w_atannode_3_w_range3262w(0) <= atannode_3_w(18);
	wire_ccc_cordic_m_w_atannode_3_w_range3270w(0) <= atannode_3_w(19);
	wire_ccc_cordic_m_w_atannode_3_w_range3126w(0) <= atannode_3_w(1);
	wire_ccc_cordic_m_w_atannode_3_w_range3278w(0) <= atannode_3_w(20);
	wire_ccc_cordic_m_w_atannode_3_w_range3286w(0) <= atannode_3_w(21);
	wire_ccc_cordic_m_w_atannode_3_w_range3294w(0) <= atannode_3_w(22);
	wire_ccc_cordic_m_w_atannode_3_w_range3302w(0) <= atannode_3_w(23);
	wire_ccc_cordic_m_w_atannode_3_w_range3310w(0) <= atannode_3_w(24);
	wire_ccc_cordic_m_w_atannode_3_w_range3318w(0) <= atannode_3_w(25);
	wire_ccc_cordic_m_w_atannode_3_w_range3326w(0) <= atannode_3_w(26);
	wire_ccc_cordic_m_w_atannode_3_w_range3334w(0) <= atannode_3_w(27);
	wire_ccc_cordic_m_w_atannode_3_w_range3342w(0) <= atannode_3_w(28);
	wire_ccc_cordic_m_w_atannode_3_w_range3350w(0) <= atannode_3_w(29);
	wire_ccc_cordic_m_w_atannode_3_w_range3134w(0) <= atannode_3_w(2);
	wire_ccc_cordic_m_w_atannode_3_w_range3358w(0) <= atannode_3_w(30);
	wire_ccc_cordic_m_w_atannode_3_w_range3366w(0) <= atannode_3_w(31);
	wire_ccc_cordic_m_w_atannode_3_w_range3374w(0) <= atannode_3_w(32);
	wire_ccc_cordic_m_w_atannode_3_w_range3382w(0) <= atannode_3_w(33);
	wire_ccc_cordic_m_w_atannode_3_w_range3142w(0) <= atannode_3_w(3);
	wire_ccc_cordic_m_w_atannode_3_w_range3150w(0) <= atannode_3_w(4);
	wire_ccc_cordic_m_w_atannode_3_w_range3158w(0) <= atannode_3_w(5);
	wire_ccc_cordic_m_w_atannode_3_w_range3166w(0) <= atannode_3_w(6);
	wire_ccc_cordic_m_w_atannode_3_w_range3174w(0) <= atannode_3_w(7);
	wire_ccc_cordic_m_w_atannode_3_w_range3182w(0) <= atannode_3_w(8);
	wire_ccc_cordic_m_w_atannode_3_w_range3190w(0) <= atannode_3_w(9);
	wire_ccc_cordic_m_w_atannode_4_w_range3954w(0) <= atannode_4_w(0);
	wire_ccc_cordic_m_w_atannode_4_w_range4035w(0) <= atannode_4_w(10);
	wire_ccc_cordic_m_w_atannode_4_w_range4043w(0) <= atannode_4_w(11);
	wire_ccc_cordic_m_w_atannode_4_w_range4051w(0) <= atannode_4_w(12);
	wire_ccc_cordic_m_w_atannode_4_w_range4059w(0) <= atannode_4_w(13);
	wire_ccc_cordic_m_w_atannode_4_w_range4067w(0) <= atannode_4_w(14);
	wire_ccc_cordic_m_w_atannode_4_w_range4075w(0) <= atannode_4_w(15);
	wire_ccc_cordic_m_w_atannode_4_w_range4083w(0) <= atannode_4_w(16);
	wire_ccc_cordic_m_w_atannode_4_w_range4091w(0) <= atannode_4_w(17);
	wire_ccc_cordic_m_w_atannode_4_w_range4099w(0) <= atannode_4_w(18);
	wire_ccc_cordic_m_w_atannode_4_w_range4107w(0) <= atannode_4_w(19);
	wire_ccc_cordic_m_w_atannode_4_w_range3963w(0) <= atannode_4_w(1);
	wire_ccc_cordic_m_w_atannode_4_w_range4115w(0) <= atannode_4_w(20);
	wire_ccc_cordic_m_w_atannode_4_w_range4123w(0) <= atannode_4_w(21);
	wire_ccc_cordic_m_w_atannode_4_w_range4131w(0) <= atannode_4_w(22);
	wire_ccc_cordic_m_w_atannode_4_w_range4139w(0) <= atannode_4_w(23);
	wire_ccc_cordic_m_w_atannode_4_w_range4147w(0) <= atannode_4_w(24);
	wire_ccc_cordic_m_w_atannode_4_w_range4155w(0) <= atannode_4_w(25);
	wire_ccc_cordic_m_w_atannode_4_w_range4163w(0) <= atannode_4_w(26);
	wire_ccc_cordic_m_w_atannode_4_w_range4171w(0) <= atannode_4_w(27);
	wire_ccc_cordic_m_w_atannode_4_w_range4179w(0) <= atannode_4_w(28);
	wire_ccc_cordic_m_w_atannode_4_w_range4187w(0) <= atannode_4_w(29);
	wire_ccc_cordic_m_w_atannode_4_w_range3971w(0) <= atannode_4_w(2);
	wire_ccc_cordic_m_w_atannode_4_w_range4195w(0) <= atannode_4_w(30);
	wire_ccc_cordic_m_w_atannode_4_w_range4203w(0) <= atannode_4_w(31);
	wire_ccc_cordic_m_w_atannode_4_w_range4211w(0) <= atannode_4_w(32);
	wire_ccc_cordic_m_w_atannode_4_w_range4219w(0) <= atannode_4_w(33);
	wire_ccc_cordic_m_w_atannode_4_w_range3979w(0) <= atannode_4_w(3);
	wire_ccc_cordic_m_w_atannode_4_w_range3987w(0) <= atannode_4_w(4);
	wire_ccc_cordic_m_w_atannode_4_w_range3995w(0) <= atannode_4_w(5);
	wire_ccc_cordic_m_w_atannode_4_w_range4003w(0) <= atannode_4_w(6);
	wire_ccc_cordic_m_w_atannode_4_w_range4011w(0) <= atannode_4_w(7);
	wire_ccc_cordic_m_w_atannode_4_w_range4019w(0) <= atannode_4_w(8);
	wire_ccc_cordic_m_w_atannode_4_w_range4027w(0) <= atannode_4_w(9);
	wire_ccc_cordic_m_w_atannode_5_w_range4786w(0) <= atannode_5_w(0);
	wire_ccc_cordic_m_w_atannode_5_w_range4867w(0) <= atannode_5_w(10);
	wire_ccc_cordic_m_w_atannode_5_w_range4875w(0) <= atannode_5_w(11);
	wire_ccc_cordic_m_w_atannode_5_w_range4883w(0) <= atannode_5_w(12);
	wire_ccc_cordic_m_w_atannode_5_w_range4891w(0) <= atannode_5_w(13);
	wire_ccc_cordic_m_w_atannode_5_w_range4899w(0) <= atannode_5_w(14);
	wire_ccc_cordic_m_w_atannode_5_w_range4907w(0) <= atannode_5_w(15);
	wire_ccc_cordic_m_w_atannode_5_w_range4915w(0) <= atannode_5_w(16);
	wire_ccc_cordic_m_w_atannode_5_w_range4923w(0) <= atannode_5_w(17);
	wire_ccc_cordic_m_w_atannode_5_w_range4931w(0) <= atannode_5_w(18);
	wire_ccc_cordic_m_w_atannode_5_w_range4939w(0) <= atannode_5_w(19);
	wire_ccc_cordic_m_w_atannode_5_w_range4795w(0) <= atannode_5_w(1);
	wire_ccc_cordic_m_w_atannode_5_w_range4947w(0) <= atannode_5_w(20);
	wire_ccc_cordic_m_w_atannode_5_w_range4955w(0) <= atannode_5_w(21);
	wire_ccc_cordic_m_w_atannode_5_w_range4963w(0) <= atannode_5_w(22);
	wire_ccc_cordic_m_w_atannode_5_w_range4971w(0) <= atannode_5_w(23);
	wire_ccc_cordic_m_w_atannode_5_w_range4979w(0) <= atannode_5_w(24);
	wire_ccc_cordic_m_w_atannode_5_w_range4987w(0) <= atannode_5_w(25);
	wire_ccc_cordic_m_w_atannode_5_w_range4995w(0) <= atannode_5_w(26);
	wire_ccc_cordic_m_w_atannode_5_w_range5003w(0) <= atannode_5_w(27);
	wire_ccc_cordic_m_w_atannode_5_w_range5011w(0) <= atannode_5_w(28);
	wire_ccc_cordic_m_w_atannode_5_w_range5019w(0) <= atannode_5_w(29);
	wire_ccc_cordic_m_w_atannode_5_w_range4803w(0) <= atannode_5_w(2);
	wire_ccc_cordic_m_w_atannode_5_w_range5027w(0) <= atannode_5_w(30);
	wire_ccc_cordic_m_w_atannode_5_w_range5035w(0) <= atannode_5_w(31);
	wire_ccc_cordic_m_w_atannode_5_w_range5043w(0) <= atannode_5_w(32);
	wire_ccc_cordic_m_w_atannode_5_w_range5051w(0) <= atannode_5_w(33);
	wire_ccc_cordic_m_w_atannode_5_w_range4811w(0) <= atannode_5_w(3);
	wire_ccc_cordic_m_w_atannode_5_w_range4819w(0) <= atannode_5_w(4);
	wire_ccc_cordic_m_w_atannode_5_w_range4827w(0) <= atannode_5_w(5);
	wire_ccc_cordic_m_w_atannode_5_w_range4835w(0) <= atannode_5_w(6);
	wire_ccc_cordic_m_w_atannode_5_w_range4843w(0) <= atannode_5_w(7);
	wire_ccc_cordic_m_w_atannode_5_w_range4851w(0) <= atannode_5_w(8);
	wire_ccc_cordic_m_w_atannode_5_w_range4859w(0) <= atannode_5_w(9);
	wire_ccc_cordic_m_w_atannode_6_w_range5613w(0) <= atannode_6_w(0);
	wire_ccc_cordic_m_w_atannode_6_w_range5694w(0) <= atannode_6_w(10);
	wire_ccc_cordic_m_w_atannode_6_w_range5702w(0) <= atannode_6_w(11);
	wire_ccc_cordic_m_w_atannode_6_w_range5710w(0) <= atannode_6_w(12);
	wire_ccc_cordic_m_w_atannode_6_w_range5718w(0) <= atannode_6_w(13);
	wire_ccc_cordic_m_w_atannode_6_w_range5726w(0) <= atannode_6_w(14);
	wire_ccc_cordic_m_w_atannode_6_w_range5734w(0) <= atannode_6_w(15);
	wire_ccc_cordic_m_w_atannode_6_w_range5742w(0) <= atannode_6_w(16);
	wire_ccc_cordic_m_w_atannode_6_w_range5750w(0) <= atannode_6_w(17);
	wire_ccc_cordic_m_w_atannode_6_w_range5758w(0) <= atannode_6_w(18);
	wire_ccc_cordic_m_w_atannode_6_w_range5766w(0) <= atannode_6_w(19);
	wire_ccc_cordic_m_w_atannode_6_w_range5622w(0) <= atannode_6_w(1);
	wire_ccc_cordic_m_w_atannode_6_w_range5774w(0) <= atannode_6_w(20);
	wire_ccc_cordic_m_w_atannode_6_w_range5782w(0) <= atannode_6_w(21);
	wire_ccc_cordic_m_w_atannode_6_w_range5790w(0) <= atannode_6_w(22);
	wire_ccc_cordic_m_w_atannode_6_w_range5798w(0) <= atannode_6_w(23);
	wire_ccc_cordic_m_w_atannode_6_w_range5806w(0) <= atannode_6_w(24);
	wire_ccc_cordic_m_w_atannode_6_w_range5814w(0) <= atannode_6_w(25);
	wire_ccc_cordic_m_w_atannode_6_w_range5822w(0) <= atannode_6_w(26);
	wire_ccc_cordic_m_w_atannode_6_w_range5830w(0) <= atannode_6_w(27);
	wire_ccc_cordic_m_w_atannode_6_w_range5838w(0) <= atannode_6_w(28);
	wire_ccc_cordic_m_w_atannode_6_w_range5846w(0) <= atannode_6_w(29);
	wire_ccc_cordic_m_w_atannode_6_w_range5630w(0) <= atannode_6_w(2);
	wire_ccc_cordic_m_w_atannode_6_w_range5854w(0) <= atannode_6_w(30);
	wire_ccc_cordic_m_w_atannode_6_w_range5862w(0) <= atannode_6_w(31);
	wire_ccc_cordic_m_w_atannode_6_w_range5870w(0) <= atannode_6_w(32);
	wire_ccc_cordic_m_w_atannode_6_w_range5878w(0) <= atannode_6_w(33);
	wire_ccc_cordic_m_w_atannode_6_w_range5638w(0) <= atannode_6_w(3);
	wire_ccc_cordic_m_w_atannode_6_w_range5646w(0) <= atannode_6_w(4);
	wire_ccc_cordic_m_w_atannode_6_w_range5654w(0) <= atannode_6_w(5);
	wire_ccc_cordic_m_w_atannode_6_w_range5662w(0) <= atannode_6_w(6);
	wire_ccc_cordic_m_w_atannode_6_w_range5670w(0) <= atannode_6_w(7);
	wire_ccc_cordic_m_w_atannode_6_w_range5678w(0) <= atannode_6_w(8);
	wire_ccc_cordic_m_w_atannode_6_w_range5686w(0) <= atannode_6_w(9);
	wire_ccc_cordic_m_w_atannode_7_w_range6435w(0) <= atannode_7_w(0);
	wire_ccc_cordic_m_w_atannode_7_w_range6516w(0) <= atannode_7_w(10);
	wire_ccc_cordic_m_w_atannode_7_w_range6524w(0) <= atannode_7_w(11);
	wire_ccc_cordic_m_w_atannode_7_w_range6532w(0) <= atannode_7_w(12);
	wire_ccc_cordic_m_w_atannode_7_w_range6540w(0) <= atannode_7_w(13);
	wire_ccc_cordic_m_w_atannode_7_w_range6548w(0) <= atannode_7_w(14);
	wire_ccc_cordic_m_w_atannode_7_w_range6556w(0) <= atannode_7_w(15);
	wire_ccc_cordic_m_w_atannode_7_w_range6564w(0) <= atannode_7_w(16);
	wire_ccc_cordic_m_w_atannode_7_w_range6572w(0) <= atannode_7_w(17);
	wire_ccc_cordic_m_w_atannode_7_w_range6580w(0) <= atannode_7_w(18);
	wire_ccc_cordic_m_w_atannode_7_w_range6588w(0) <= atannode_7_w(19);
	wire_ccc_cordic_m_w_atannode_7_w_range6444w(0) <= atannode_7_w(1);
	wire_ccc_cordic_m_w_atannode_7_w_range6596w(0) <= atannode_7_w(20);
	wire_ccc_cordic_m_w_atannode_7_w_range6604w(0) <= atannode_7_w(21);
	wire_ccc_cordic_m_w_atannode_7_w_range6612w(0) <= atannode_7_w(22);
	wire_ccc_cordic_m_w_atannode_7_w_range6620w(0) <= atannode_7_w(23);
	wire_ccc_cordic_m_w_atannode_7_w_range6628w(0) <= atannode_7_w(24);
	wire_ccc_cordic_m_w_atannode_7_w_range6636w(0) <= atannode_7_w(25);
	wire_ccc_cordic_m_w_atannode_7_w_range6644w(0) <= atannode_7_w(26);
	wire_ccc_cordic_m_w_atannode_7_w_range6652w(0) <= atannode_7_w(27);
	wire_ccc_cordic_m_w_atannode_7_w_range6660w(0) <= atannode_7_w(28);
	wire_ccc_cordic_m_w_atannode_7_w_range6668w(0) <= atannode_7_w(29);
	wire_ccc_cordic_m_w_atannode_7_w_range6452w(0) <= atannode_7_w(2);
	wire_ccc_cordic_m_w_atannode_7_w_range6676w(0) <= atannode_7_w(30);
	wire_ccc_cordic_m_w_atannode_7_w_range6684w(0) <= atannode_7_w(31);
	wire_ccc_cordic_m_w_atannode_7_w_range6692w(0) <= atannode_7_w(32);
	wire_ccc_cordic_m_w_atannode_7_w_range6700w(0) <= atannode_7_w(33);
	wire_ccc_cordic_m_w_atannode_7_w_range6460w(0) <= atannode_7_w(3);
	wire_ccc_cordic_m_w_atannode_7_w_range6468w(0) <= atannode_7_w(4);
	wire_ccc_cordic_m_w_atannode_7_w_range6476w(0) <= atannode_7_w(5);
	wire_ccc_cordic_m_w_atannode_7_w_range6484w(0) <= atannode_7_w(6);
	wire_ccc_cordic_m_w_atannode_7_w_range6492w(0) <= atannode_7_w(7);
	wire_ccc_cordic_m_w_atannode_7_w_range6500w(0) <= atannode_7_w(8);
	wire_ccc_cordic_m_w_atannode_7_w_range6508w(0) <= atannode_7_w(9);
	wire_ccc_cordic_m_w_atannode_8_w_range7252w(0) <= atannode_8_w(0);
	wire_ccc_cordic_m_w_atannode_8_w_range7333w(0) <= atannode_8_w(10);
	wire_ccc_cordic_m_w_atannode_8_w_range7341w(0) <= atannode_8_w(11);
	wire_ccc_cordic_m_w_atannode_8_w_range7349w(0) <= atannode_8_w(12);
	wire_ccc_cordic_m_w_atannode_8_w_range7357w(0) <= atannode_8_w(13);
	wire_ccc_cordic_m_w_atannode_8_w_range7365w(0) <= atannode_8_w(14);
	wire_ccc_cordic_m_w_atannode_8_w_range7373w(0) <= atannode_8_w(15);
	wire_ccc_cordic_m_w_atannode_8_w_range7381w(0) <= atannode_8_w(16);
	wire_ccc_cordic_m_w_atannode_8_w_range7389w(0) <= atannode_8_w(17);
	wire_ccc_cordic_m_w_atannode_8_w_range7397w(0) <= atannode_8_w(18);
	wire_ccc_cordic_m_w_atannode_8_w_range7405w(0) <= atannode_8_w(19);
	wire_ccc_cordic_m_w_atannode_8_w_range7261w(0) <= atannode_8_w(1);
	wire_ccc_cordic_m_w_atannode_8_w_range7413w(0) <= atannode_8_w(20);
	wire_ccc_cordic_m_w_atannode_8_w_range7421w(0) <= atannode_8_w(21);
	wire_ccc_cordic_m_w_atannode_8_w_range7429w(0) <= atannode_8_w(22);
	wire_ccc_cordic_m_w_atannode_8_w_range7437w(0) <= atannode_8_w(23);
	wire_ccc_cordic_m_w_atannode_8_w_range7445w(0) <= atannode_8_w(24);
	wire_ccc_cordic_m_w_atannode_8_w_range7453w(0) <= atannode_8_w(25);
	wire_ccc_cordic_m_w_atannode_8_w_range7461w(0) <= atannode_8_w(26);
	wire_ccc_cordic_m_w_atannode_8_w_range7469w(0) <= atannode_8_w(27);
	wire_ccc_cordic_m_w_atannode_8_w_range7477w(0) <= atannode_8_w(28);
	wire_ccc_cordic_m_w_atannode_8_w_range7485w(0) <= atannode_8_w(29);
	wire_ccc_cordic_m_w_atannode_8_w_range7269w(0) <= atannode_8_w(2);
	wire_ccc_cordic_m_w_atannode_8_w_range7493w(0) <= atannode_8_w(30);
	wire_ccc_cordic_m_w_atannode_8_w_range7501w(0) <= atannode_8_w(31);
	wire_ccc_cordic_m_w_atannode_8_w_range7509w(0) <= atannode_8_w(32);
	wire_ccc_cordic_m_w_atannode_8_w_range7517w(0) <= atannode_8_w(33);
	wire_ccc_cordic_m_w_atannode_8_w_range7277w(0) <= atannode_8_w(3);
	wire_ccc_cordic_m_w_atannode_8_w_range7285w(0) <= atannode_8_w(4);
	wire_ccc_cordic_m_w_atannode_8_w_range7293w(0) <= atannode_8_w(5);
	wire_ccc_cordic_m_w_atannode_8_w_range7301w(0) <= atannode_8_w(6);
	wire_ccc_cordic_m_w_atannode_8_w_range7309w(0) <= atannode_8_w(7);
	wire_ccc_cordic_m_w_atannode_8_w_range7317w(0) <= atannode_8_w(8);
	wire_ccc_cordic_m_w_atannode_8_w_range7325w(0) <= atannode_8_w(9);
	wire_ccc_cordic_m_w_atannode_9_w_range8064w(0) <= atannode_9_w(0);
	wire_ccc_cordic_m_w_atannode_9_w_range8145w(0) <= atannode_9_w(10);
	wire_ccc_cordic_m_w_atannode_9_w_range8153w(0) <= atannode_9_w(11);
	wire_ccc_cordic_m_w_atannode_9_w_range8161w(0) <= atannode_9_w(12);
	wire_ccc_cordic_m_w_atannode_9_w_range8169w(0) <= atannode_9_w(13);
	wire_ccc_cordic_m_w_atannode_9_w_range8177w(0) <= atannode_9_w(14);
	wire_ccc_cordic_m_w_atannode_9_w_range8185w(0) <= atannode_9_w(15);
	wire_ccc_cordic_m_w_atannode_9_w_range8193w(0) <= atannode_9_w(16);
	wire_ccc_cordic_m_w_atannode_9_w_range8201w(0) <= atannode_9_w(17);
	wire_ccc_cordic_m_w_atannode_9_w_range8209w(0) <= atannode_9_w(18);
	wire_ccc_cordic_m_w_atannode_9_w_range8217w(0) <= atannode_9_w(19);
	wire_ccc_cordic_m_w_atannode_9_w_range8073w(0) <= atannode_9_w(1);
	wire_ccc_cordic_m_w_atannode_9_w_range8225w(0) <= atannode_9_w(20);
	wire_ccc_cordic_m_w_atannode_9_w_range8233w(0) <= atannode_9_w(21);
	wire_ccc_cordic_m_w_atannode_9_w_range8241w(0) <= atannode_9_w(22);
	wire_ccc_cordic_m_w_atannode_9_w_range8249w(0) <= atannode_9_w(23);
	wire_ccc_cordic_m_w_atannode_9_w_range8257w(0) <= atannode_9_w(24);
	wire_ccc_cordic_m_w_atannode_9_w_range8265w(0) <= atannode_9_w(25);
	wire_ccc_cordic_m_w_atannode_9_w_range8273w(0) <= atannode_9_w(26);
	wire_ccc_cordic_m_w_atannode_9_w_range8281w(0) <= atannode_9_w(27);
	wire_ccc_cordic_m_w_atannode_9_w_range8289w(0) <= atannode_9_w(28);
	wire_ccc_cordic_m_w_atannode_9_w_range8297w(0) <= atannode_9_w(29);
	wire_ccc_cordic_m_w_atannode_9_w_range8081w(0) <= atannode_9_w(2);
	wire_ccc_cordic_m_w_atannode_9_w_range8305w(0) <= atannode_9_w(30);
	wire_ccc_cordic_m_w_atannode_9_w_range8313w(0) <= atannode_9_w(31);
	wire_ccc_cordic_m_w_atannode_9_w_range8321w(0) <= atannode_9_w(32);
	wire_ccc_cordic_m_w_atannode_9_w_range8329w(0) <= atannode_9_w(33);
	wire_ccc_cordic_m_w_atannode_9_w_range8089w(0) <= atannode_9_w(3);
	wire_ccc_cordic_m_w_atannode_9_w_range8097w(0) <= atannode_9_w(4);
	wire_ccc_cordic_m_w_atannode_9_w_range8105w(0) <= atannode_9_w(5);
	wire_ccc_cordic_m_w_atannode_9_w_range8113w(0) <= atannode_9_w(6);
	wire_ccc_cordic_m_w_atannode_9_w_range8121w(0) <= atannode_9_w(7);
	wire_ccc_cordic_m_w_atannode_9_w_range8129w(0) <= atannode_9_w(8);
	wire_ccc_cordic_m_w_atannode_9_w_range8137w(0) <= atannode_9_w(9);
	wire_ccc_cordic_m_w_pre_estimate_w_range10751w(0) <= pre_estimate_w(0);
	wire_ccc_cordic_m_w_pre_estimate_w_range10794w(0) <= pre_estimate_w(10);
	wire_ccc_cordic_m_w_pre_estimate_w_range10799w(0) <= pre_estimate_w(11);
	wire_ccc_cordic_m_w_pre_estimate_w_range10804w(0) <= pre_estimate_w(12);
	wire_ccc_cordic_m_w_pre_estimate_w_range10809w(0) <= pre_estimate_w(13);
	wire_ccc_cordic_m_w_pre_estimate_w_range10814w(0) <= pre_estimate_w(14);
	wire_ccc_cordic_m_w_pre_estimate_w_range10819w(0) <= pre_estimate_w(15);
	wire_ccc_cordic_m_w_pre_estimate_w_range10824w(0) <= pre_estimate_w(16);
	wire_ccc_cordic_m_w_pre_estimate_w_range10829w(0) <= pre_estimate_w(17);
	wire_ccc_cordic_m_w_pre_estimate_w_range10834w(0) <= pre_estimate_w(18);
	wire_ccc_cordic_m_w_pre_estimate_w_range10839w(0) <= pre_estimate_w(19);
	wire_ccc_cordic_m_w_pre_estimate_w_range10759w(0) <= pre_estimate_w(1);
	wire_ccc_cordic_m_w_pre_estimate_w_range10844w(0) <= pre_estimate_w(20);
	wire_ccc_cordic_m_w_pre_estimate_w_range10849w(0) <= pre_estimate_w(21);
	wire_ccc_cordic_m_w_pre_estimate_w_range10854w(0) <= pre_estimate_w(22);
	wire_ccc_cordic_m_w_pre_estimate_w_range10859w(0) <= pre_estimate_w(23);
	wire_ccc_cordic_m_w_pre_estimate_w_range10864w(0) <= pre_estimate_w(24);
	wire_ccc_cordic_m_w_pre_estimate_w_range10869w(0) <= pre_estimate_w(25);
	wire_ccc_cordic_m_w_pre_estimate_w_range10874w(0) <= pre_estimate_w(26);
	wire_ccc_cordic_m_w_pre_estimate_w_range10879w(0) <= pre_estimate_w(27);
	wire_ccc_cordic_m_w_pre_estimate_w_range10884w(0) <= pre_estimate_w(28);
	wire_ccc_cordic_m_w_pre_estimate_w_range10889w(0) <= pre_estimate_w(29);
	wire_ccc_cordic_m_w_pre_estimate_w_range10750w(0) <= pre_estimate_w(2);
	wire_ccc_cordic_m_w_pre_estimate_w_range10894w(0) <= pre_estimate_w(30);
	wire_ccc_cordic_m_w_pre_estimate_w_range10899w(0) <= pre_estimate_w(31);
	wire_ccc_cordic_m_w_pre_estimate_w_range10904w(0) <= pre_estimate_w(32);
	wire_ccc_cordic_m_w_pre_estimate_w_range10909w(0) <= pre_estimate_w(33);
	wire_ccc_cordic_m_w_pre_estimate_w_range10758w(0) <= pre_estimate_w(3);
	wire_ccc_cordic_m_w_pre_estimate_w_range10764w(0) <= pre_estimate_w(4);
	wire_ccc_cordic_m_w_pre_estimate_w_range10769w(0) <= pre_estimate_w(5);
	wire_ccc_cordic_m_w_pre_estimate_w_range10774w(0) <= pre_estimate_w(6);
	wire_ccc_cordic_m_w_pre_estimate_w_range10779w(0) <= pre_estimate_w(7);
	wire_ccc_cordic_m_w_pre_estimate_w_range10784w(0) <= pre_estimate_w(8);
	wire_ccc_cordic_m_w_pre_estimate_w_range10789w(0) <= pre_estimate_w(9);
	wire_ccc_cordic_m_w_radians_range410w(0) <= radians(0);
	wire_ccc_cordic_m_w_radians_range458w(0) <= radians(10);
	wire_ccc_cordic_m_w_radians_range463w(0) <= radians(11);
	wire_ccc_cordic_m_w_radians_range468w(0) <= radians(12);
	wire_ccc_cordic_m_w_radians_range473w(0) <= radians(13);
	wire_ccc_cordic_m_w_radians_range478w(0) <= radians(14);
	wire_ccc_cordic_m_w_radians_range483w(0) <= radians(15);
	wire_ccc_cordic_m_w_radians_range488w(0) <= radians(16);
	wire_ccc_cordic_m_w_radians_range493w(0) <= radians(17);
	wire_ccc_cordic_m_w_radians_range498w(0) <= radians(18);
	wire_ccc_cordic_m_w_radians_range503w(0) <= radians(19);
	wire_ccc_cordic_m_w_radians_range415w(0) <= radians(1);
	wire_ccc_cordic_m_w_radians_range508w(0) <= radians(20);
	wire_ccc_cordic_m_w_radians_range513w(0) <= radians(21);
	wire_ccc_cordic_m_w_radians_range518w(0) <= radians(22);
	wire_ccc_cordic_m_w_radians_range523w(0) <= radians(23);
	wire_ccc_cordic_m_w_radians_range528w(0) <= radians(24);
	wire_ccc_cordic_m_w_radians_range533w(0) <= radians(25);
	wire_ccc_cordic_m_w_radians_range538w(0) <= radians(26);
	wire_ccc_cordic_m_w_radians_range543w(0) <= radians(27);
	wire_ccc_cordic_m_w_radians_range548w(0) <= radians(28);
	wire_ccc_cordic_m_w_radians_range553w(0) <= radians(29);
	wire_ccc_cordic_m_w_radians_range418w(0) <= radians(2);
	wire_ccc_cordic_m_w_radians_range558w(0) <= radians(30);
	wire_ccc_cordic_m_w_radians_range563w(0) <= radians(31);
	wire_ccc_cordic_m_w_radians_range568w(0) <= radians(32);
	wire_ccc_cordic_m_w_radians_range573w(0) <= radians(33);
	wire_ccc_cordic_m_w_radians_range423w(0) <= radians(3);
	wire_ccc_cordic_m_w_radians_range428w(0) <= radians(4);
	wire_ccc_cordic_m_w_radians_range433w(0) <= radians(5);
	wire_ccc_cordic_m_w_radians_range438w(0) <= radians(6);
	wire_ccc_cordic_m_w_radians_range443w(0) <= radians(7);
	wire_ccc_cordic_m_w_radians_range448w(0) <= radians(8);
	wire_ccc_cordic_m_w_radians_range453w(0) <= radians(9);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7782w(0) <= x_prenode_10_w(0);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7865w(0) <= x_prenode_10_w(10);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7873w(0) <= x_prenode_10_w(11);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7881w(0) <= x_prenode_10_w(12);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7889w(0) <= x_prenode_10_w(13);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7897w(0) <= x_prenode_10_w(14);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7905w(0) <= x_prenode_10_w(15);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7913w(0) <= x_prenode_10_w(16);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7921w(0) <= x_prenode_10_w(17);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7929w(0) <= x_prenode_10_w(18);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7937w(0) <= x_prenode_10_w(19);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7793w(0) <= x_prenode_10_w(1);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7945w(0) <= x_prenode_10_w(20);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7953w(0) <= x_prenode_10_w(21);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7961w(0) <= x_prenode_10_w(22);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7969w(0) <= x_prenode_10_w(23);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7977w(0) <= x_prenode_10_w(24);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7985w(0) <= x_prenode_10_w(25);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7993w(0) <= x_prenode_10_w(26);
	wire_ccc_cordic_m_w_x_prenode_10_w_range8001w(0) <= x_prenode_10_w(27);
	wire_ccc_cordic_m_w_x_prenode_10_w_range8009w(0) <= x_prenode_10_w(28);
	wire_ccc_cordic_m_w_x_prenode_10_w_range8017w(0) <= x_prenode_10_w(29);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7801w(0) <= x_prenode_10_w(2);
	wire_ccc_cordic_m_w_x_prenode_10_w_range8025w(0) <= x_prenode_10_w(30);
	wire_ccc_cordic_m_w_x_prenode_10_w_range8033w(0) <= x_prenode_10_w(31);
	wire_ccc_cordic_m_w_x_prenode_10_w_range8041w(0) <= x_prenode_10_w(32);
	wire_ccc_cordic_m_w_x_prenode_10_w_range8049w(0) <= x_prenode_10_w(33);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7809w(0) <= x_prenode_10_w(3);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7817w(0) <= x_prenode_10_w(4);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7825w(0) <= x_prenode_10_w(5);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7833w(0) <= x_prenode_10_w(6);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7841w(0) <= x_prenode_10_w(7);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7849w(0) <= x_prenode_10_w(8);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7857w(0) <= x_prenode_10_w(9);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8589w(0) <= x_prenode_11_w(0);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8672w(0) <= x_prenode_11_w(10);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8680w(0) <= x_prenode_11_w(11);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8688w(0) <= x_prenode_11_w(12);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8696w(0) <= x_prenode_11_w(13);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8704w(0) <= x_prenode_11_w(14);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8712w(0) <= x_prenode_11_w(15);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8720w(0) <= x_prenode_11_w(16);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8728w(0) <= x_prenode_11_w(17);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8736w(0) <= x_prenode_11_w(18);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8744w(0) <= x_prenode_11_w(19);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8600w(0) <= x_prenode_11_w(1);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8752w(0) <= x_prenode_11_w(20);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8760w(0) <= x_prenode_11_w(21);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8768w(0) <= x_prenode_11_w(22);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8776w(0) <= x_prenode_11_w(23);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8784w(0) <= x_prenode_11_w(24);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8792w(0) <= x_prenode_11_w(25);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8800w(0) <= x_prenode_11_w(26);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8808w(0) <= x_prenode_11_w(27);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8816w(0) <= x_prenode_11_w(28);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8824w(0) <= x_prenode_11_w(29);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8608w(0) <= x_prenode_11_w(2);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8832w(0) <= x_prenode_11_w(30);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8840w(0) <= x_prenode_11_w(31);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8848w(0) <= x_prenode_11_w(32);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8856w(0) <= x_prenode_11_w(33);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8616w(0) <= x_prenode_11_w(3);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8624w(0) <= x_prenode_11_w(4);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8632w(0) <= x_prenode_11_w(5);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8640w(0) <= x_prenode_11_w(6);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8648w(0) <= x_prenode_11_w(7);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8656w(0) <= x_prenode_11_w(8);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8664w(0) <= x_prenode_11_w(9);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9391w(0) <= x_prenode_12_w(0);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9474w(0) <= x_prenode_12_w(10);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9482w(0) <= x_prenode_12_w(11);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9490w(0) <= x_prenode_12_w(12);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9498w(0) <= x_prenode_12_w(13);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9506w(0) <= x_prenode_12_w(14);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9514w(0) <= x_prenode_12_w(15);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9522w(0) <= x_prenode_12_w(16);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9530w(0) <= x_prenode_12_w(17);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9538w(0) <= x_prenode_12_w(18);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9546w(0) <= x_prenode_12_w(19);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9402w(0) <= x_prenode_12_w(1);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9554w(0) <= x_prenode_12_w(20);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9562w(0) <= x_prenode_12_w(21);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9570w(0) <= x_prenode_12_w(22);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9578w(0) <= x_prenode_12_w(23);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9586w(0) <= x_prenode_12_w(24);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9594w(0) <= x_prenode_12_w(25);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9602w(0) <= x_prenode_12_w(26);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9610w(0) <= x_prenode_12_w(27);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9618w(0) <= x_prenode_12_w(28);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9626w(0) <= x_prenode_12_w(29);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9410w(0) <= x_prenode_12_w(2);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9634w(0) <= x_prenode_12_w(30);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9642w(0) <= x_prenode_12_w(31);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9650w(0) <= x_prenode_12_w(32);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9658w(0) <= x_prenode_12_w(33);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9418w(0) <= x_prenode_12_w(3);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9426w(0) <= x_prenode_12_w(4);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9434w(0) <= x_prenode_12_w(5);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9442w(0) <= x_prenode_12_w(6);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9450w(0) <= x_prenode_12_w(7);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9458w(0) <= x_prenode_12_w(8);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9466w(0) <= x_prenode_12_w(9);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10188w(0) <= x_prenode_13_w(0);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10271w(0) <= x_prenode_13_w(10);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10279w(0) <= x_prenode_13_w(11);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10287w(0) <= x_prenode_13_w(12);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10295w(0) <= x_prenode_13_w(13);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10303w(0) <= x_prenode_13_w(14);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10311w(0) <= x_prenode_13_w(15);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10319w(0) <= x_prenode_13_w(16);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10327w(0) <= x_prenode_13_w(17);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10335w(0) <= x_prenode_13_w(18);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10343w(0) <= x_prenode_13_w(19);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10199w(0) <= x_prenode_13_w(1);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10351w(0) <= x_prenode_13_w(20);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10359w(0) <= x_prenode_13_w(21);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10367w(0) <= x_prenode_13_w(22);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10375w(0) <= x_prenode_13_w(23);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10383w(0) <= x_prenode_13_w(24);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10391w(0) <= x_prenode_13_w(25);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10399w(0) <= x_prenode_13_w(26);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10407w(0) <= x_prenode_13_w(27);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10415w(0) <= x_prenode_13_w(28);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10423w(0) <= x_prenode_13_w(29);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10207w(0) <= x_prenode_13_w(2);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10431w(0) <= x_prenode_13_w(30);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10439w(0) <= x_prenode_13_w(31);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10447w(0) <= x_prenode_13_w(32);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10455w(0) <= x_prenode_13_w(33);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10215w(0) <= x_prenode_13_w(3);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10223w(0) <= x_prenode_13_w(4);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10231w(0) <= x_prenode_13_w(5);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10239w(0) <= x_prenode_13_w(6);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10247w(0) <= x_prenode_13_w(7);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10255w(0) <= x_prenode_13_w(8);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10263w(0) <= x_prenode_13_w(9);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1146w(0) <= x_prenode_2_w(0);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1229w(0) <= x_prenode_2_w(10);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1237w(0) <= x_prenode_2_w(11);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1245w(0) <= x_prenode_2_w(12);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1253w(0) <= x_prenode_2_w(13);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1261w(0) <= x_prenode_2_w(14);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1269w(0) <= x_prenode_2_w(15);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1277w(0) <= x_prenode_2_w(16);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1285w(0) <= x_prenode_2_w(17);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1293w(0) <= x_prenode_2_w(18);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1301w(0) <= x_prenode_2_w(19);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1157w(0) <= x_prenode_2_w(1);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1309w(0) <= x_prenode_2_w(20);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1317w(0) <= x_prenode_2_w(21);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1325w(0) <= x_prenode_2_w(22);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1333w(0) <= x_prenode_2_w(23);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1341w(0) <= x_prenode_2_w(24);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1349w(0) <= x_prenode_2_w(25);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1357w(0) <= x_prenode_2_w(26);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1365w(0) <= x_prenode_2_w(27);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1373w(0) <= x_prenode_2_w(28);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1381w(0) <= x_prenode_2_w(29);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1165w(0) <= x_prenode_2_w(2);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1389w(0) <= x_prenode_2_w(30);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1397w(0) <= x_prenode_2_w(31);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1405w(0) <= x_prenode_2_w(32);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1413w(0) <= x_prenode_2_w(33);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1173w(0) <= x_prenode_2_w(3);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1181w(0) <= x_prenode_2_w(4);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1189w(0) <= x_prenode_2_w(5);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1197w(0) <= x_prenode_2_w(6);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1205w(0) <= x_prenode_2_w(7);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1213w(0) <= x_prenode_2_w(8);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1221w(0) <= x_prenode_2_w(9);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1993w(0) <= x_prenode_3_w(0);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2076w(0) <= x_prenode_3_w(10);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2084w(0) <= x_prenode_3_w(11);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2092w(0) <= x_prenode_3_w(12);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2100w(0) <= x_prenode_3_w(13);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2108w(0) <= x_prenode_3_w(14);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2116w(0) <= x_prenode_3_w(15);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2124w(0) <= x_prenode_3_w(16);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2132w(0) <= x_prenode_3_w(17);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2140w(0) <= x_prenode_3_w(18);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2148w(0) <= x_prenode_3_w(19);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2004w(0) <= x_prenode_3_w(1);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2156w(0) <= x_prenode_3_w(20);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2164w(0) <= x_prenode_3_w(21);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2172w(0) <= x_prenode_3_w(22);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2180w(0) <= x_prenode_3_w(23);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2188w(0) <= x_prenode_3_w(24);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2196w(0) <= x_prenode_3_w(25);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2204w(0) <= x_prenode_3_w(26);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2212w(0) <= x_prenode_3_w(27);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2220w(0) <= x_prenode_3_w(28);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2228w(0) <= x_prenode_3_w(29);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2012w(0) <= x_prenode_3_w(2);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2236w(0) <= x_prenode_3_w(30);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2244w(0) <= x_prenode_3_w(31);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2252w(0) <= x_prenode_3_w(32);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2260w(0) <= x_prenode_3_w(33);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2020w(0) <= x_prenode_3_w(3);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2028w(0) <= x_prenode_3_w(4);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2036w(0) <= x_prenode_3_w(5);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2044w(0) <= x_prenode_3_w(6);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2052w(0) <= x_prenode_3_w(7);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2060w(0) <= x_prenode_3_w(8);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2068w(0) <= x_prenode_3_w(9);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2835w(0) <= x_prenode_4_w(0);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2918w(0) <= x_prenode_4_w(10);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2926w(0) <= x_prenode_4_w(11);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2934w(0) <= x_prenode_4_w(12);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2942w(0) <= x_prenode_4_w(13);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2950w(0) <= x_prenode_4_w(14);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2958w(0) <= x_prenode_4_w(15);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2966w(0) <= x_prenode_4_w(16);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2974w(0) <= x_prenode_4_w(17);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2982w(0) <= x_prenode_4_w(18);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2990w(0) <= x_prenode_4_w(19);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2846w(0) <= x_prenode_4_w(1);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2998w(0) <= x_prenode_4_w(20);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3006w(0) <= x_prenode_4_w(21);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3014w(0) <= x_prenode_4_w(22);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3022w(0) <= x_prenode_4_w(23);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3030w(0) <= x_prenode_4_w(24);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3038w(0) <= x_prenode_4_w(25);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3046w(0) <= x_prenode_4_w(26);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3054w(0) <= x_prenode_4_w(27);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3062w(0) <= x_prenode_4_w(28);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3070w(0) <= x_prenode_4_w(29);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2854w(0) <= x_prenode_4_w(2);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3078w(0) <= x_prenode_4_w(30);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3086w(0) <= x_prenode_4_w(31);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3094w(0) <= x_prenode_4_w(32);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3102w(0) <= x_prenode_4_w(33);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2862w(0) <= x_prenode_4_w(3);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2870w(0) <= x_prenode_4_w(4);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2878w(0) <= x_prenode_4_w(5);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2886w(0) <= x_prenode_4_w(6);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2894w(0) <= x_prenode_4_w(7);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2902w(0) <= x_prenode_4_w(8);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2910w(0) <= x_prenode_4_w(9);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3672w(0) <= x_prenode_5_w(0);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3755w(0) <= x_prenode_5_w(10);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3763w(0) <= x_prenode_5_w(11);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3771w(0) <= x_prenode_5_w(12);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3779w(0) <= x_prenode_5_w(13);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3787w(0) <= x_prenode_5_w(14);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3795w(0) <= x_prenode_5_w(15);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3803w(0) <= x_prenode_5_w(16);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3811w(0) <= x_prenode_5_w(17);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3819w(0) <= x_prenode_5_w(18);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3827w(0) <= x_prenode_5_w(19);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3683w(0) <= x_prenode_5_w(1);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3835w(0) <= x_prenode_5_w(20);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3843w(0) <= x_prenode_5_w(21);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3851w(0) <= x_prenode_5_w(22);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3859w(0) <= x_prenode_5_w(23);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3867w(0) <= x_prenode_5_w(24);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3875w(0) <= x_prenode_5_w(25);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3883w(0) <= x_prenode_5_w(26);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3891w(0) <= x_prenode_5_w(27);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3899w(0) <= x_prenode_5_w(28);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3907w(0) <= x_prenode_5_w(29);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3691w(0) <= x_prenode_5_w(2);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3915w(0) <= x_prenode_5_w(30);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3923w(0) <= x_prenode_5_w(31);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3931w(0) <= x_prenode_5_w(32);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3939w(0) <= x_prenode_5_w(33);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3699w(0) <= x_prenode_5_w(3);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3707w(0) <= x_prenode_5_w(4);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3715w(0) <= x_prenode_5_w(5);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3723w(0) <= x_prenode_5_w(6);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3731w(0) <= x_prenode_5_w(7);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3739w(0) <= x_prenode_5_w(8);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3747w(0) <= x_prenode_5_w(9);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4504w(0) <= x_prenode_6_w(0);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4587w(0) <= x_prenode_6_w(10);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4595w(0) <= x_prenode_6_w(11);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4603w(0) <= x_prenode_6_w(12);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4611w(0) <= x_prenode_6_w(13);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4619w(0) <= x_prenode_6_w(14);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4627w(0) <= x_prenode_6_w(15);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4635w(0) <= x_prenode_6_w(16);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4643w(0) <= x_prenode_6_w(17);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4651w(0) <= x_prenode_6_w(18);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4659w(0) <= x_prenode_6_w(19);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4515w(0) <= x_prenode_6_w(1);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4667w(0) <= x_prenode_6_w(20);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4675w(0) <= x_prenode_6_w(21);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4683w(0) <= x_prenode_6_w(22);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4691w(0) <= x_prenode_6_w(23);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4699w(0) <= x_prenode_6_w(24);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4707w(0) <= x_prenode_6_w(25);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4715w(0) <= x_prenode_6_w(26);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4723w(0) <= x_prenode_6_w(27);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4731w(0) <= x_prenode_6_w(28);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4739w(0) <= x_prenode_6_w(29);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4523w(0) <= x_prenode_6_w(2);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4747w(0) <= x_prenode_6_w(30);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4755w(0) <= x_prenode_6_w(31);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4763w(0) <= x_prenode_6_w(32);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4771w(0) <= x_prenode_6_w(33);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4531w(0) <= x_prenode_6_w(3);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4539w(0) <= x_prenode_6_w(4);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4547w(0) <= x_prenode_6_w(5);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4555w(0) <= x_prenode_6_w(6);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4563w(0) <= x_prenode_6_w(7);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4571w(0) <= x_prenode_6_w(8);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4579w(0) <= x_prenode_6_w(9);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5331w(0) <= x_prenode_7_w(0);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5414w(0) <= x_prenode_7_w(10);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5422w(0) <= x_prenode_7_w(11);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5430w(0) <= x_prenode_7_w(12);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5438w(0) <= x_prenode_7_w(13);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5446w(0) <= x_prenode_7_w(14);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5454w(0) <= x_prenode_7_w(15);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5462w(0) <= x_prenode_7_w(16);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5470w(0) <= x_prenode_7_w(17);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5478w(0) <= x_prenode_7_w(18);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5486w(0) <= x_prenode_7_w(19);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5342w(0) <= x_prenode_7_w(1);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5494w(0) <= x_prenode_7_w(20);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5502w(0) <= x_prenode_7_w(21);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5510w(0) <= x_prenode_7_w(22);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5518w(0) <= x_prenode_7_w(23);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5526w(0) <= x_prenode_7_w(24);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5534w(0) <= x_prenode_7_w(25);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5542w(0) <= x_prenode_7_w(26);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5550w(0) <= x_prenode_7_w(27);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5558w(0) <= x_prenode_7_w(28);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5566w(0) <= x_prenode_7_w(29);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5350w(0) <= x_prenode_7_w(2);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5574w(0) <= x_prenode_7_w(30);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5582w(0) <= x_prenode_7_w(31);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5590w(0) <= x_prenode_7_w(32);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5598w(0) <= x_prenode_7_w(33);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5358w(0) <= x_prenode_7_w(3);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5366w(0) <= x_prenode_7_w(4);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5374w(0) <= x_prenode_7_w(5);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5382w(0) <= x_prenode_7_w(6);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5390w(0) <= x_prenode_7_w(7);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5398w(0) <= x_prenode_7_w(8);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5406w(0) <= x_prenode_7_w(9);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6153w(0) <= x_prenode_8_w(0);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6236w(0) <= x_prenode_8_w(10);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6244w(0) <= x_prenode_8_w(11);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6252w(0) <= x_prenode_8_w(12);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6260w(0) <= x_prenode_8_w(13);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6268w(0) <= x_prenode_8_w(14);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6276w(0) <= x_prenode_8_w(15);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6284w(0) <= x_prenode_8_w(16);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6292w(0) <= x_prenode_8_w(17);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6300w(0) <= x_prenode_8_w(18);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6308w(0) <= x_prenode_8_w(19);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6164w(0) <= x_prenode_8_w(1);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6316w(0) <= x_prenode_8_w(20);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6324w(0) <= x_prenode_8_w(21);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6332w(0) <= x_prenode_8_w(22);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6340w(0) <= x_prenode_8_w(23);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6348w(0) <= x_prenode_8_w(24);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6356w(0) <= x_prenode_8_w(25);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6364w(0) <= x_prenode_8_w(26);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6372w(0) <= x_prenode_8_w(27);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6380w(0) <= x_prenode_8_w(28);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6388w(0) <= x_prenode_8_w(29);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6172w(0) <= x_prenode_8_w(2);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6396w(0) <= x_prenode_8_w(30);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6404w(0) <= x_prenode_8_w(31);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6412w(0) <= x_prenode_8_w(32);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6420w(0) <= x_prenode_8_w(33);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6180w(0) <= x_prenode_8_w(3);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6188w(0) <= x_prenode_8_w(4);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6196w(0) <= x_prenode_8_w(5);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6204w(0) <= x_prenode_8_w(6);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6212w(0) <= x_prenode_8_w(7);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6220w(0) <= x_prenode_8_w(8);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6228w(0) <= x_prenode_8_w(9);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6970w(0) <= x_prenode_9_w(0);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7053w(0) <= x_prenode_9_w(10);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7061w(0) <= x_prenode_9_w(11);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7069w(0) <= x_prenode_9_w(12);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7077w(0) <= x_prenode_9_w(13);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7085w(0) <= x_prenode_9_w(14);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7093w(0) <= x_prenode_9_w(15);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7101w(0) <= x_prenode_9_w(16);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7109w(0) <= x_prenode_9_w(17);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7117w(0) <= x_prenode_9_w(18);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7125w(0) <= x_prenode_9_w(19);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6981w(0) <= x_prenode_9_w(1);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7133w(0) <= x_prenode_9_w(20);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7141w(0) <= x_prenode_9_w(21);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7149w(0) <= x_prenode_9_w(22);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7157w(0) <= x_prenode_9_w(23);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7165w(0) <= x_prenode_9_w(24);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7173w(0) <= x_prenode_9_w(25);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7181w(0) <= x_prenode_9_w(26);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7189w(0) <= x_prenode_9_w(27);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7197w(0) <= x_prenode_9_w(28);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7205w(0) <= x_prenode_9_w(29);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6989w(0) <= x_prenode_9_w(2);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7213w(0) <= x_prenode_9_w(30);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7221w(0) <= x_prenode_9_w(31);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7229w(0) <= x_prenode_9_w(32);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7237w(0) <= x_prenode_9_w(33);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6997w(0) <= x_prenode_9_w(3);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7005w(0) <= x_prenode_9_w(4);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7013w(0) <= x_prenode_9_w(5);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7021w(0) <= x_prenode_9_w(6);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7029w(0) <= x_prenode_9_w(7);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7037w(0) <= x_prenode_9_w(8);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7045w(0) <= x_prenode_9_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7569w(0) <= x_prenodeone_10_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7628w(0) <= x_prenodeone_10_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7634w(0) <= x_prenodeone_10_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7640w(0) <= x_prenodeone_10_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7646w(0) <= x_prenodeone_10_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7652w(0) <= x_prenodeone_10_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7658w(0) <= x_prenodeone_10_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7664w(0) <= x_prenodeone_10_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7670w(0) <= x_prenodeone_10_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7676w(0) <= x_prenodeone_10_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7682w(0) <= x_prenodeone_10_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7574w(0) <= x_prenodeone_10_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7688w(0) <= x_prenodeone_10_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7694w(0) <= x_prenodeone_10_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7700w(0) <= x_prenodeone_10_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7706w(0) <= x_prenodeone_10_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7711w(0) <= x_prenodeone_10_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7522w(0) <= x_prenodeone_10_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7528w(0) <= x_prenodeone_10_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7530w(0) <= x_prenodeone_10_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7532w(0) <= x_prenodeone_10_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7534w(0) <= x_prenodeone_10_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7580w(0) <= x_prenodeone_10_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7536w(0) <= x_prenodeone_10_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7538w(0) <= x_prenodeone_10_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7540w(0) <= x_prenodeone_10_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7542w(0) <= x_prenodeone_10_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7586w(0) <= x_prenodeone_10_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7592w(0) <= x_prenodeone_10_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7598w(0) <= x_prenodeone_10_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7604w(0) <= x_prenodeone_10_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7610w(0) <= x_prenodeone_10_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7616w(0) <= x_prenodeone_10_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7622w(0) <= x_prenodeone_10_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8385w(0) <= x_prenodeone_11_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8444w(0) <= x_prenodeone_11_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8450w(0) <= x_prenodeone_11_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8456w(0) <= x_prenodeone_11_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8462w(0) <= x_prenodeone_11_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8468w(0) <= x_prenodeone_11_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8474w(0) <= x_prenodeone_11_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8480w(0) <= x_prenodeone_11_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8486w(0) <= x_prenodeone_11_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8492w(0) <= x_prenodeone_11_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8498w(0) <= x_prenodeone_11_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8390w(0) <= x_prenodeone_11_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8504w(0) <= x_prenodeone_11_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8510w(0) <= x_prenodeone_11_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8516w(0) <= x_prenodeone_11_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8521w(0) <= x_prenodeone_11_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8334w(0) <= x_prenodeone_11_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8340w(0) <= x_prenodeone_11_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8342w(0) <= x_prenodeone_11_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8344w(0) <= x_prenodeone_11_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8346w(0) <= x_prenodeone_11_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8348w(0) <= x_prenodeone_11_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8396w(0) <= x_prenodeone_11_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8350w(0) <= x_prenodeone_11_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8352w(0) <= x_prenodeone_11_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8354w(0) <= x_prenodeone_11_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8356w(0) <= x_prenodeone_11_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8402w(0) <= x_prenodeone_11_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8408w(0) <= x_prenodeone_11_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8414w(0) <= x_prenodeone_11_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8420w(0) <= x_prenodeone_11_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8426w(0) <= x_prenodeone_11_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8432w(0) <= x_prenodeone_11_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8438w(0) <= x_prenodeone_11_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9196w(0) <= x_prenodeone_12_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9255w(0) <= x_prenodeone_12_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9261w(0) <= x_prenodeone_12_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9267w(0) <= x_prenodeone_12_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9273w(0) <= x_prenodeone_12_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9279w(0) <= x_prenodeone_12_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9285w(0) <= x_prenodeone_12_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9291w(0) <= x_prenodeone_12_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9297w(0) <= x_prenodeone_12_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9303w(0) <= x_prenodeone_12_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9309w(0) <= x_prenodeone_12_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9201w(0) <= x_prenodeone_12_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9315w(0) <= x_prenodeone_12_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9321w(0) <= x_prenodeone_12_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9326w(0) <= x_prenodeone_12_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9141w(0) <= x_prenodeone_12_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9147w(0) <= x_prenodeone_12_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9149w(0) <= x_prenodeone_12_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9151w(0) <= x_prenodeone_12_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9153w(0) <= x_prenodeone_12_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9155w(0) <= x_prenodeone_12_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9157w(0) <= x_prenodeone_12_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9207w(0) <= x_prenodeone_12_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9159w(0) <= x_prenodeone_12_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9161w(0) <= x_prenodeone_12_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9163w(0) <= x_prenodeone_12_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9165w(0) <= x_prenodeone_12_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9213w(0) <= x_prenodeone_12_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9219w(0) <= x_prenodeone_12_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9225w(0) <= x_prenodeone_12_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9231w(0) <= x_prenodeone_12_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9237w(0) <= x_prenodeone_12_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9243w(0) <= x_prenodeone_12_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9249w(0) <= x_prenodeone_12_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10002w(0) <= x_prenodeone_13_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10061w(0) <= x_prenodeone_13_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10067w(0) <= x_prenodeone_13_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10073w(0) <= x_prenodeone_13_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10079w(0) <= x_prenodeone_13_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10085w(0) <= x_prenodeone_13_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10091w(0) <= x_prenodeone_13_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10097w(0) <= x_prenodeone_13_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10103w(0) <= x_prenodeone_13_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10109w(0) <= x_prenodeone_13_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10115w(0) <= x_prenodeone_13_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10007w(0) <= x_prenodeone_13_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10121w(0) <= x_prenodeone_13_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10126w(0) <= x_prenodeone_13_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9943w(0) <= x_prenodeone_13_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9949w(0) <= x_prenodeone_13_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9951w(0) <= x_prenodeone_13_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9953w(0) <= x_prenodeone_13_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9955w(0) <= x_prenodeone_13_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9957w(0) <= x_prenodeone_13_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9959w(0) <= x_prenodeone_13_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9961w(0) <= x_prenodeone_13_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10013w(0) <= x_prenodeone_13_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9963w(0) <= x_prenodeone_13_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9965w(0) <= x_prenodeone_13_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9967w(0) <= x_prenodeone_13_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9969w(0) <= x_prenodeone_13_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10019w(0) <= x_prenodeone_13_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10025w(0) <= x_prenodeone_13_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10031w(0) <= x_prenodeone_13_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10037w(0) <= x_prenodeone_13_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10043w(0) <= x_prenodeone_13_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10049w(0) <= x_prenodeone_13_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10055w(0) <= x_prenodeone_13_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range861w(0) <= x_prenodeone_2_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range920w(0) <= x_prenodeone_2_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range926w(0) <= x_prenodeone_2_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range932w(0) <= x_prenodeone_2_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range938w(0) <= x_prenodeone_2_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range944w(0) <= x_prenodeone_2_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range950w(0) <= x_prenodeone_2_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range956w(0) <= x_prenodeone_2_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range962w(0) <= x_prenodeone_2_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range968w(0) <= x_prenodeone_2_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range974w(0) <= x_prenodeone_2_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range866w(0) <= x_prenodeone_2_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range980w(0) <= x_prenodeone_2_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range986w(0) <= x_prenodeone_2_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range992w(0) <= x_prenodeone_2_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range998w(0) <= x_prenodeone_2_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range1004w(0) <= x_prenodeone_2_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range1010w(0) <= x_prenodeone_2_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range1016w(0) <= x_prenodeone_2_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range1022w(0) <= x_prenodeone_2_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range1028w(0) <= x_prenodeone_2_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range1034w(0) <= x_prenodeone_2_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range872w(0) <= x_prenodeone_2_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range1040w(0) <= x_prenodeone_2_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range1046w(0) <= x_prenodeone_2_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range1051w(0) <= x_prenodeone_2_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range846w(0) <= x_prenodeone_2_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range878w(0) <= x_prenodeone_2_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range884w(0) <= x_prenodeone_2_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range890w(0) <= x_prenodeone_2_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range896w(0) <= x_prenodeone_2_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range902w(0) <= x_prenodeone_2_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range908w(0) <= x_prenodeone_2_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range914w(0) <= x_prenodeone_2_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1717w(0) <= x_prenodeone_3_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1776w(0) <= x_prenodeone_3_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1782w(0) <= x_prenodeone_3_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1788w(0) <= x_prenodeone_3_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1794w(0) <= x_prenodeone_3_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1800w(0) <= x_prenodeone_3_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1806w(0) <= x_prenodeone_3_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1812w(0) <= x_prenodeone_3_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1818w(0) <= x_prenodeone_3_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1824w(0) <= x_prenodeone_3_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1830w(0) <= x_prenodeone_3_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1722w(0) <= x_prenodeone_3_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1836w(0) <= x_prenodeone_3_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1842w(0) <= x_prenodeone_3_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1848w(0) <= x_prenodeone_3_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1854w(0) <= x_prenodeone_3_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1860w(0) <= x_prenodeone_3_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1866w(0) <= x_prenodeone_3_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1872w(0) <= x_prenodeone_3_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1878w(0) <= x_prenodeone_3_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1884w(0) <= x_prenodeone_3_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1890w(0) <= x_prenodeone_3_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1728w(0) <= x_prenodeone_3_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1896w(0) <= x_prenodeone_3_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1901w(0) <= x_prenodeone_3_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1698w(0) <= x_prenodeone_3_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1704w(0) <= x_prenodeone_3_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1734w(0) <= x_prenodeone_3_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1740w(0) <= x_prenodeone_3_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1746w(0) <= x_prenodeone_3_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1752w(0) <= x_prenodeone_3_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1758w(0) <= x_prenodeone_3_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1764w(0) <= x_prenodeone_3_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1770w(0) <= x_prenodeone_3_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2568w(0) <= x_prenodeone_4_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2627w(0) <= x_prenodeone_4_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2633w(0) <= x_prenodeone_4_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2639w(0) <= x_prenodeone_4_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2645w(0) <= x_prenodeone_4_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2651w(0) <= x_prenodeone_4_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2657w(0) <= x_prenodeone_4_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2663w(0) <= x_prenodeone_4_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2669w(0) <= x_prenodeone_4_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2675w(0) <= x_prenodeone_4_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2681w(0) <= x_prenodeone_4_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2573w(0) <= x_prenodeone_4_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2687w(0) <= x_prenodeone_4_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2693w(0) <= x_prenodeone_4_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2699w(0) <= x_prenodeone_4_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2705w(0) <= x_prenodeone_4_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2711w(0) <= x_prenodeone_4_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2717w(0) <= x_prenodeone_4_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2723w(0) <= x_prenodeone_4_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2729w(0) <= x_prenodeone_4_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2735w(0) <= x_prenodeone_4_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2741w(0) <= x_prenodeone_4_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2579w(0) <= x_prenodeone_4_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2746w(0) <= x_prenodeone_4_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2545w(0) <= x_prenodeone_4_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2551w(0) <= x_prenodeone_4_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2553w(0) <= x_prenodeone_4_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2585w(0) <= x_prenodeone_4_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2591w(0) <= x_prenodeone_4_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2597w(0) <= x_prenodeone_4_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2603w(0) <= x_prenodeone_4_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2609w(0) <= x_prenodeone_4_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2615w(0) <= x_prenodeone_4_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2621w(0) <= x_prenodeone_4_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3414w(0) <= x_prenodeone_5_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3473w(0) <= x_prenodeone_5_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3479w(0) <= x_prenodeone_5_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3485w(0) <= x_prenodeone_5_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3491w(0) <= x_prenodeone_5_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3497w(0) <= x_prenodeone_5_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3503w(0) <= x_prenodeone_5_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3509w(0) <= x_prenodeone_5_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3515w(0) <= x_prenodeone_5_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3521w(0) <= x_prenodeone_5_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3527w(0) <= x_prenodeone_5_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3419w(0) <= x_prenodeone_5_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3533w(0) <= x_prenodeone_5_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3539w(0) <= x_prenodeone_5_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3545w(0) <= x_prenodeone_5_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3551w(0) <= x_prenodeone_5_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3557w(0) <= x_prenodeone_5_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3563w(0) <= x_prenodeone_5_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3569w(0) <= x_prenodeone_5_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3575w(0) <= x_prenodeone_5_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3581w(0) <= x_prenodeone_5_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3586w(0) <= x_prenodeone_5_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3425w(0) <= x_prenodeone_5_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3387w(0) <= x_prenodeone_5_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3393w(0) <= x_prenodeone_5_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3395w(0) <= x_prenodeone_5_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3397w(0) <= x_prenodeone_5_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3431w(0) <= x_prenodeone_5_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3437w(0) <= x_prenodeone_5_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3443w(0) <= x_prenodeone_5_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3449w(0) <= x_prenodeone_5_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3455w(0) <= x_prenodeone_5_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3461w(0) <= x_prenodeone_5_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3467w(0) <= x_prenodeone_5_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4255w(0) <= x_prenodeone_6_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4314w(0) <= x_prenodeone_6_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4320w(0) <= x_prenodeone_6_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4326w(0) <= x_prenodeone_6_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4332w(0) <= x_prenodeone_6_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4338w(0) <= x_prenodeone_6_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4344w(0) <= x_prenodeone_6_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4350w(0) <= x_prenodeone_6_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4356w(0) <= x_prenodeone_6_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4362w(0) <= x_prenodeone_6_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4368w(0) <= x_prenodeone_6_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4260w(0) <= x_prenodeone_6_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4374w(0) <= x_prenodeone_6_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4380w(0) <= x_prenodeone_6_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4386w(0) <= x_prenodeone_6_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4392w(0) <= x_prenodeone_6_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4398w(0) <= x_prenodeone_6_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4404w(0) <= x_prenodeone_6_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4410w(0) <= x_prenodeone_6_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4416w(0) <= x_prenodeone_6_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4421w(0) <= x_prenodeone_6_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4224w(0) <= x_prenodeone_6_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4266w(0) <= x_prenodeone_6_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4230w(0) <= x_prenodeone_6_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4232w(0) <= x_prenodeone_6_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4234w(0) <= x_prenodeone_6_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4236w(0) <= x_prenodeone_6_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4272w(0) <= x_prenodeone_6_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4278w(0) <= x_prenodeone_6_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4284w(0) <= x_prenodeone_6_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4290w(0) <= x_prenodeone_6_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4296w(0) <= x_prenodeone_6_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4302w(0) <= x_prenodeone_6_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4308w(0) <= x_prenodeone_6_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5091w(0) <= x_prenodeone_7_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5150w(0) <= x_prenodeone_7_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5156w(0) <= x_prenodeone_7_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5162w(0) <= x_prenodeone_7_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5168w(0) <= x_prenodeone_7_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5174w(0) <= x_prenodeone_7_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5180w(0) <= x_prenodeone_7_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5186w(0) <= x_prenodeone_7_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5192w(0) <= x_prenodeone_7_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5198w(0) <= x_prenodeone_7_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5204w(0) <= x_prenodeone_7_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5096w(0) <= x_prenodeone_7_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5210w(0) <= x_prenodeone_7_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5216w(0) <= x_prenodeone_7_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5222w(0) <= x_prenodeone_7_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5228w(0) <= x_prenodeone_7_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5234w(0) <= x_prenodeone_7_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5240w(0) <= x_prenodeone_7_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5246w(0) <= x_prenodeone_7_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5251w(0) <= x_prenodeone_7_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5056w(0) <= x_prenodeone_7_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5062w(0) <= x_prenodeone_7_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5102w(0) <= x_prenodeone_7_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5064w(0) <= x_prenodeone_7_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5066w(0) <= x_prenodeone_7_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5068w(0) <= x_prenodeone_7_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5070w(0) <= x_prenodeone_7_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5108w(0) <= x_prenodeone_7_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5114w(0) <= x_prenodeone_7_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5120w(0) <= x_prenodeone_7_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5126w(0) <= x_prenodeone_7_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5132w(0) <= x_prenodeone_7_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5138w(0) <= x_prenodeone_7_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5144w(0) <= x_prenodeone_7_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5922w(0) <= x_prenodeone_8_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5981w(0) <= x_prenodeone_8_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5987w(0) <= x_prenodeone_8_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5993w(0) <= x_prenodeone_8_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5999w(0) <= x_prenodeone_8_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6005w(0) <= x_prenodeone_8_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6011w(0) <= x_prenodeone_8_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6017w(0) <= x_prenodeone_8_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6023w(0) <= x_prenodeone_8_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6029w(0) <= x_prenodeone_8_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6035w(0) <= x_prenodeone_8_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5927w(0) <= x_prenodeone_8_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6041w(0) <= x_prenodeone_8_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6047w(0) <= x_prenodeone_8_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6053w(0) <= x_prenodeone_8_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6059w(0) <= x_prenodeone_8_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6065w(0) <= x_prenodeone_8_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6071w(0) <= x_prenodeone_8_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6076w(0) <= x_prenodeone_8_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5883w(0) <= x_prenodeone_8_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5889w(0) <= x_prenodeone_8_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5891w(0) <= x_prenodeone_8_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5933w(0) <= x_prenodeone_8_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5893w(0) <= x_prenodeone_8_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5895w(0) <= x_prenodeone_8_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5897w(0) <= x_prenodeone_8_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5899w(0) <= x_prenodeone_8_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5939w(0) <= x_prenodeone_8_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5945w(0) <= x_prenodeone_8_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5951w(0) <= x_prenodeone_8_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5957w(0) <= x_prenodeone_8_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5963w(0) <= x_prenodeone_8_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5969w(0) <= x_prenodeone_8_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5975w(0) <= x_prenodeone_8_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6748w(0) <= x_prenodeone_9_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6807w(0) <= x_prenodeone_9_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6813w(0) <= x_prenodeone_9_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6819w(0) <= x_prenodeone_9_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6825w(0) <= x_prenodeone_9_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6831w(0) <= x_prenodeone_9_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6837w(0) <= x_prenodeone_9_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6843w(0) <= x_prenodeone_9_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6849w(0) <= x_prenodeone_9_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6855w(0) <= x_prenodeone_9_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6861w(0) <= x_prenodeone_9_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6753w(0) <= x_prenodeone_9_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6867w(0) <= x_prenodeone_9_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6873w(0) <= x_prenodeone_9_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6879w(0) <= x_prenodeone_9_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6885w(0) <= x_prenodeone_9_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6891w(0) <= x_prenodeone_9_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6896w(0) <= x_prenodeone_9_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6705w(0) <= x_prenodeone_9_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6711w(0) <= x_prenodeone_9_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6713w(0) <= x_prenodeone_9_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6715w(0) <= x_prenodeone_9_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6759w(0) <= x_prenodeone_9_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6717w(0) <= x_prenodeone_9_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6719w(0) <= x_prenodeone_9_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6721w(0) <= x_prenodeone_9_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6723w(0) <= x_prenodeone_9_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6765w(0) <= x_prenodeone_9_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6771w(0) <= x_prenodeone_9_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6777w(0) <= x_prenodeone_9_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6783w(0) <= x_prenodeone_9_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6789w(0) <= x_prenodeone_9_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6795w(0) <= x_prenodeone_9_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6801w(0) <= x_prenodeone_9_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7714w(0) <= x_prenodetwo_10_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7743w(0) <= x_prenodetwo_10_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7746w(0) <= x_prenodetwo_10_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7749w(0) <= x_prenodetwo_10_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7752w(0) <= x_prenodetwo_10_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7755w(0) <= x_prenodetwo_10_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7758w(0) <= x_prenodetwo_10_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7761w(0) <= x_prenodetwo_10_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7764w(0) <= x_prenodetwo_10_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7767w(0) <= x_prenodetwo_10_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7770w(0) <= x_prenodetwo_10_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7716w(0) <= x_prenodetwo_10_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7773w(0) <= x_prenodetwo_10_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7776w(0) <= x_prenodetwo_10_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7779w(0) <= x_prenodetwo_10_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7544w(0) <= x_prenodetwo_10_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7548w(0) <= x_prenodetwo_10_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7550w(0) <= x_prenodetwo_10_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7552w(0) <= x_prenodetwo_10_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7554w(0) <= x_prenodetwo_10_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7556w(0) <= x_prenodetwo_10_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7558w(0) <= x_prenodetwo_10_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7719w(0) <= x_prenodetwo_10_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7560w(0) <= x_prenodetwo_10_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7562w(0) <= x_prenodetwo_10_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7564w(0) <= x_prenodetwo_10_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7566w(0) <= x_prenodetwo_10_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7722w(0) <= x_prenodetwo_10_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7725w(0) <= x_prenodetwo_10_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7728w(0) <= x_prenodetwo_10_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7731w(0) <= x_prenodetwo_10_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7734w(0) <= x_prenodetwo_10_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7737w(0) <= x_prenodetwo_10_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7740w(0) <= x_prenodetwo_10_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8524w(0) <= x_prenodetwo_11_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8553w(0) <= x_prenodetwo_11_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8556w(0) <= x_prenodetwo_11_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8559w(0) <= x_prenodetwo_11_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8562w(0) <= x_prenodetwo_11_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8565w(0) <= x_prenodetwo_11_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8568w(0) <= x_prenodetwo_11_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8571w(0) <= x_prenodetwo_11_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8574w(0) <= x_prenodetwo_11_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8577w(0) <= x_prenodetwo_11_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8580w(0) <= x_prenodetwo_11_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8526w(0) <= x_prenodetwo_11_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8583w(0) <= x_prenodetwo_11_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8586w(0) <= x_prenodetwo_11_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8358w(0) <= x_prenodetwo_11_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8362w(0) <= x_prenodetwo_11_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8364w(0) <= x_prenodetwo_11_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8366w(0) <= x_prenodetwo_11_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8368w(0) <= x_prenodetwo_11_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8370w(0) <= x_prenodetwo_11_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8372w(0) <= x_prenodetwo_11_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8374w(0) <= x_prenodetwo_11_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8529w(0) <= x_prenodetwo_11_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8376w(0) <= x_prenodetwo_11_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8378w(0) <= x_prenodetwo_11_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8380w(0) <= x_prenodetwo_11_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8382w(0) <= x_prenodetwo_11_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8532w(0) <= x_prenodetwo_11_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8535w(0) <= x_prenodetwo_11_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8538w(0) <= x_prenodetwo_11_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8541w(0) <= x_prenodetwo_11_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8544w(0) <= x_prenodetwo_11_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8547w(0) <= x_prenodetwo_11_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8550w(0) <= x_prenodetwo_11_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9329w(0) <= x_prenodetwo_12_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9358w(0) <= x_prenodetwo_12_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9361w(0) <= x_prenodetwo_12_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9364w(0) <= x_prenodetwo_12_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9367w(0) <= x_prenodetwo_12_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9370w(0) <= x_prenodetwo_12_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9373w(0) <= x_prenodetwo_12_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9376w(0) <= x_prenodetwo_12_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9379w(0) <= x_prenodetwo_12_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9382w(0) <= x_prenodetwo_12_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9385w(0) <= x_prenodetwo_12_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9331w(0) <= x_prenodetwo_12_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9388w(0) <= x_prenodetwo_12_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9167w(0) <= x_prenodetwo_12_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9171w(0) <= x_prenodetwo_12_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9173w(0) <= x_prenodetwo_12_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9175w(0) <= x_prenodetwo_12_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9177w(0) <= x_prenodetwo_12_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9179w(0) <= x_prenodetwo_12_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9181w(0) <= x_prenodetwo_12_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9183w(0) <= x_prenodetwo_12_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9185w(0) <= x_prenodetwo_12_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9334w(0) <= x_prenodetwo_12_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9187w(0) <= x_prenodetwo_12_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9189w(0) <= x_prenodetwo_12_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9191w(0) <= x_prenodetwo_12_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9193w(0) <= x_prenodetwo_12_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9337w(0) <= x_prenodetwo_12_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9340w(0) <= x_prenodetwo_12_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9343w(0) <= x_prenodetwo_12_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9346w(0) <= x_prenodetwo_12_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9349w(0) <= x_prenodetwo_12_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9352w(0) <= x_prenodetwo_12_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9355w(0) <= x_prenodetwo_12_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10129w(0) <= x_prenodetwo_13_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10158w(0) <= x_prenodetwo_13_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10161w(0) <= x_prenodetwo_13_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10164w(0) <= x_prenodetwo_13_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10167w(0) <= x_prenodetwo_13_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10170w(0) <= x_prenodetwo_13_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10173w(0) <= x_prenodetwo_13_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10176w(0) <= x_prenodetwo_13_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10179w(0) <= x_prenodetwo_13_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10182w(0) <= x_prenodetwo_13_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10185w(0) <= x_prenodetwo_13_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10131w(0) <= x_prenodetwo_13_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9971w(0) <= x_prenodetwo_13_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9975w(0) <= x_prenodetwo_13_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9977w(0) <= x_prenodetwo_13_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9979w(0) <= x_prenodetwo_13_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9981w(0) <= x_prenodetwo_13_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9983w(0) <= x_prenodetwo_13_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9985w(0) <= x_prenodetwo_13_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9987w(0) <= x_prenodetwo_13_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9989w(0) <= x_prenodetwo_13_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9991w(0) <= x_prenodetwo_13_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10134w(0) <= x_prenodetwo_13_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9993w(0) <= x_prenodetwo_13_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9995w(0) <= x_prenodetwo_13_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9997w(0) <= x_prenodetwo_13_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9999w(0) <= x_prenodetwo_13_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10137w(0) <= x_prenodetwo_13_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10140w(0) <= x_prenodetwo_13_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10143w(0) <= x_prenodetwo_13_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10146w(0) <= x_prenodetwo_13_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10149w(0) <= x_prenodetwo_13_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10152w(0) <= x_prenodetwo_13_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10155w(0) <= x_prenodetwo_13_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1054w(0) <= x_prenodetwo_2_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1083w(0) <= x_prenodetwo_2_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1086w(0) <= x_prenodetwo_2_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1089w(0) <= x_prenodetwo_2_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1092w(0) <= x_prenodetwo_2_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1095w(0) <= x_prenodetwo_2_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1098w(0) <= x_prenodetwo_2_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1101w(0) <= x_prenodetwo_2_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1104w(0) <= x_prenodetwo_2_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1107w(0) <= x_prenodetwo_2_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1110w(0) <= x_prenodetwo_2_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1056w(0) <= x_prenodetwo_2_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1113w(0) <= x_prenodetwo_2_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1116w(0) <= x_prenodetwo_2_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1119w(0) <= x_prenodetwo_2_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1122w(0) <= x_prenodetwo_2_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1125w(0) <= x_prenodetwo_2_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1128w(0) <= x_prenodetwo_2_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1131w(0) <= x_prenodetwo_2_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1134w(0) <= x_prenodetwo_2_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1137w(0) <= x_prenodetwo_2_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1140w(0) <= x_prenodetwo_2_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1059w(0) <= x_prenodetwo_2_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1143w(0) <= x_prenodetwo_2_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range852w(0) <= x_prenodetwo_2_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range856w(0) <= x_prenodetwo_2_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range858w(0) <= x_prenodetwo_2_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1062w(0) <= x_prenodetwo_2_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1065w(0) <= x_prenodetwo_2_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1068w(0) <= x_prenodetwo_2_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1071w(0) <= x_prenodetwo_2_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1074w(0) <= x_prenodetwo_2_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1077w(0) <= x_prenodetwo_2_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1080w(0) <= x_prenodetwo_2_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1904w(0) <= x_prenodetwo_3_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1933w(0) <= x_prenodetwo_3_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1936w(0) <= x_prenodetwo_3_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1939w(0) <= x_prenodetwo_3_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1942w(0) <= x_prenodetwo_3_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1945w(0) <= x_prenodetwo_3_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1948w(0) <= x_prenodetwo_3_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1951w(0) <= x_prenodetwo_3_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1954w(0) <= x_prenodetwo_3_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1957w(0) <= x_prenodetwo_3_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1960w(0) <= x_prenodetwo_3_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1906w(0) <= x_prenodetwo_3_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1963w(0) <= x_prenodetwo_3_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1966w(0) <= x_prenodetwo_3_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1969w(0) <= x_prenodetwo_3_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1972w(0) <= x_prenodetwo_3_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1975w(0) <= x_prenodetwo_3_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1978w(0) <= x_prenodetwo_3_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1981w(0) <= x_prenodetwo_3_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1984w(0) <= x_prenodetwo_3_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1987w(0) <= x_prenodetwo_3_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1990w(0) <= x_prenodetwo_3_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1909w(0) <= x_prenodetwo_3_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1706w(0) <= x_prenodetwo_3_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1710w(0) <= x_prenodetwo_3_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1712w(0) <= x_prenodetwo_3_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1714w(0) <= x_prenodetwo_3_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1912w(0) <= x_prenodetwo_3_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1915w(0) <= x_prenodetwo_3_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1918w(0) <= x_prenodetwo_3_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1921w(0) <= x_prenodetwo_3_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1924w(0) <= x_prenodetwo_3_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1927w(0) <= x_prenodetwo_3_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1930w(0) <= x_prenodetwo_3_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2749w(0) <= x_prenodetwo_4_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2778w(0) <= x_prenodetwo_4_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2781w(0) <= x_prenodetwo_4_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2784w(0) <= x_prenodetwo_4_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2787w(0) <= x_prenodetwo_4_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2790w(0) <= x_prenodetwo_4_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2793w(0) <= x_prenodetwo_4_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2796w(0) <= x_prenodetwo_4_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2799w(0) <= x_prenodetwo_4_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2802w(0) <= x_prenodetwo_4_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2805w(0) <= x_prenodetwo_4_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2751w(0) <= x_prenodetwo_4_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2808w(0) <= x_prenodetwo_4_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2811w(0) <= x_prenodetwo_4_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2814w(0) <= x_prenodetwo_4_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2817w(0) <= x_prenodetwo_4_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2820w(0) <= x_prenodetwo_4_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2823w(0) <= x_prenodetwo_4_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2826w(0) <= x_prenodetwo_4_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2829w(0) <= x_prenodetwo_4_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2832w(0) <= x_prenodetwo_4_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2555w(0) <= x_prenodetwo_4_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2754w(0) <= x_prenodetwo_4_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2559w(0) <= x_prenodetwo_4_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2561w(0) <= x_prenodetwo_4_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2563w(0) <= x_prenodetwo_4_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2565w(0) <= x_prenodetwo_4_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2757w(0) <= x_prenodetwo_4_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2760w(0) <= x_prenodetwo_4_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2763w(0) <= x_prenodetwo_4_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2766w(0) <= x_prenodetwo_4_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2769w(0) <= x_prenodetwo_4_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2772w(0) <= x_prenodetwo_4_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2775w(0) <= x_prenodetwo_4_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3589w(0) <= x_prenodetwo_5_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3618w(0) <= x_prenodetwo_5_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3621w(0) <= x_prenodetwo_5_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3624w(0) <= x_prenodetwo_5_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3627w(0) <= x_prenodetwo_5_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3630w(0) <= x_prenodetwo_5_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3633w(0) <= x_prenodetwo_5_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3636w(0) <= x_prenodetwo_5_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3639w(0) <= x_prenodetwo_5_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3642w(0) <= x_prenodetwo_5_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3645w(0) <= x_prenodetwo_5_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3591w(0) <= x_prenodetwo_5_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3648w(0) <= x_prenodetwo_5_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3651w(0) <= x_prenodetwo_5_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3654w(0) <= x_prenodetwo_5_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3657w(0) <= x_prenodetwo_5_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3660w(0) <= x_prenodetwo_5_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3663w(0) <= x_prenodetwo_5_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3666w(0) <= x_prenodetwo_5_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3669w(0) <= x_prenodetwo_5_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3399w(0) <= x_prenodetwo_5_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3403w(0) <= x_prenodetwo_5_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3594w(0) <= x_prenodetwo_5_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3405w(0) <= x_prenodetwo_5_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3407w(0) <= x_prenodetwo_5_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3409w(0) <= x_prenodetwo_5_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3411w(0) <= x_prenodetwo_5_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3597w(0) <= x_prenodetwo_5_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3600w(0) <= x_prenodetwo_5_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3603w(0) <= x_prenodetwo_5_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3606w(0) <= x_prenodetwo_5_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3609w(0) <= x_prenodetwo_5_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3612w(0) <= x_prenodetwo_5_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3615w(0) <= x_prenodetwo_5_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4424w(0) <= x_prenodetwo_6_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4453w(0) <= x_prenodetwo_6_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4456w(0) <= x_prenodetwo_6_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4459w(0) <= x_prenodetwo_6_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4462w(0) <= x_prenodetwo_6_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4465w(0) <= x_prenodetwo_6_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4468w(0) <= x_prenodetwo_6_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4471w(0) <= x_prenodetwo_6_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4474w(0) <= x_prenodetwo_6_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4477w(0) <= x_prenodetwo_6_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4480w(0) <= x_prenodetwo_6_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4426w(0) <= x_prenodetwo_6_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4483w(0) <= x_prenodetwo_6_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4486w(0) <= x_prenodetwo_6_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4489w(0) <= x_prenodetwo_6_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4492w(0) <= x_prenodetwo_6_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4495w(0) <= x_prenodetwo_6_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4498w(0) <= x_prenodetwo_6_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4501w(0) <= x_prenodetwo_6_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4238w(0) <= x_prenodetwo_6_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4242w(0) <= x_prenodetwo_6_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4244w(0) <= x_prenodetwo_6_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4429w(0) <= x_prenodetwo_6_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4246w(0) <= x_prenodetwo_6_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4248w(0) <= x_prenodetwo_6_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4250w(0) <= x_prenodetwo_6_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4252w(0) <= x_prenodetwo_6_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4432w(0) <= x_prenodetwo_6_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4435w(0) <= x_prenodetwo_6_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4438w(0) <= x_prenodetwo_6_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4441w(0) <= x_prenodetwo_6_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4444w(0) <= x_prenodetwo_6_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4447w(0) <= x_prenodetwo_6_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4450w(0) <= x_prenodetwo_6_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5254w(0) <= x_prenodetwo_7_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5283w(0) <= x_prenodetwo_7_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5286w(0) <= x_prenodetwo_7_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5289w(0) <= x_prenodetwo_7_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5292w(0) <= x_prenodetwo_7_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5295w(0) <= x_prenodetwo_7_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5298w(0) <= x_prenodetwo_7_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5301w(0) <= x_prenodetwo_7_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5304w(0) <= x_prenodetwo_7_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5307w(0) <= x_prenodetwo_7_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5310w(0) <= x_prenodetwo_7_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5256w(0) <= x_prenodetwo_7_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5313w(0) <= x_prenodetwo_7_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5316w(0) <= x_prenodetwo_7_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5319w(0) <= x_prenodetwo_7_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5322w(0) <= x_prenodetwo_7_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5325w(0) <= x_prenodetwo_7_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5328w(0) <= x_prenodetwo_7_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5072w(0) <= x_prenodetwo_7_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5076w(0) <= x_prenodetwo_7_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5078w(0) <= x_prenodetwo_7_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5080w(0) <= x_prenodetwo_7_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5259w(0) <= x_prenodetwo_7_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5082w(0) <= x_prenodetwo_7_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5084w(0) <= x_prenodetwo_7_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5086w(0) <= x_prenodetwo_7_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5088w(0) <= x_prenodetwo_7_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5262w(0) <= x_prenodetwo_7_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5265w(0) <= x_prenodetwo_7_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5268w(0) <= x_prenodetwo_7_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5271w(0) <= x_prenodetwo_7_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5274w(0) <= x_prenodetwo_7_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5277w(0) <= x_prenodetwo_7_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5280w(0) <= x_prenodetwo_7_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6079w(0) <= x_prenodetwo_8_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6108w(0) <= x_prenodetwo_8_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6111w(0) <= x_prenodetwo_8_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6114w(0) <= x_prenodetwo_8_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6117w(0) <= x_prenodetwo_8_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6120w(0) <= x_prenodetwo_8_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6123w(0) <= x_prenodetwo_8_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6126w(0) <= x_prenodetwo_8_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6129w(0) <= x_prenodetwo_8_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6132w(0) <= x_prenodetwo_8_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6135w(0) <= x_prenodetwo_8_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6081w(0) <= x_prenodetwo_8_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6138w(0) <= x_prenodetwo_8_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6141w(0) <= x_prenodetwo_8_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6144w(0) <= x_prenodetwo_8_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6147w(0) <= x_prenodetwo_8_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6150w(0) <= x_prenodetwo_8_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5901w(0) <= x_prenodetwo_8_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5905w(0) <= x_prenodetwo_8_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5907w(0) <= x_prenodetwo_8_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5909w(0) <= x_prenodetwo_8_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5911w(0) <= x_prenodetwo_8_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6084w(0) <= x_prenodetwo_8_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5913w(0) <= x_prenodetwo_8_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5915w(0) <= x_prenodetwo_8_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5917w(0) <= x_prenodetwo_8_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5919w(0) <= x_prenodetwo_8_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6087w(0) <= x_prenodetwo_8_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6090w(0) <= x_prenodetwo_8_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6093w(0) <= x_prenodetwo_8_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6096w(0) <= x_prenodetwo_8_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6099w(0) <= x_prenodetwo_8_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6102w(0) <= x_prenodetwo_8_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6105w(0) <= x_prenodetwo_8_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6899w(0) <= x_prenodetwo_9_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6928w(0) <= x_prenodetwo_9_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6931w(0) <= x_prenodetwo_9_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6934w(0) <= x_prenodetwo_9_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6937w(0) <= x_prenodetwo_9_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6940w(0) <= x_prenodetwo_9_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6943w(0) <= x_prenodetwo_9_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6946w(0) <= x_prenodetwo_9_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6949w(0) <= x_prenodetwo_9_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6952w(0) <= x_prenodetwo_9_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6955w(0) <= x_prenodetwo_9_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6901w(0) <= x_prenodetwo_9_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6958w(0) <= x_prenodetwo_9_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6961w(0) <= x_prenodetwo_9_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6964w(0) <= x_prenodetwo_9_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6967w(0) <= x_prenodetwo_9_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6725w(0) <= x_prenodetwo_9_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6729w(0) <= x_prenodetwo_9_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6731w(0) <= x_prenodetwo_9_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6733w(0) <= x_prenodetwo_9_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6735w(0) <= x_prenodetwo_9_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6737w(0) <= x_prenodetwo_9_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6904w(0) <= x_prenodetwo_9_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6739w(0) <= x_prenodetwo_9_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6741w(0) <= x_prenodetwo_9_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6743w(0) <= x_prenodetwo_9_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6745w(0) <= x_prenodetwo_9_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6907w(0) <= x_prenodetwo_9_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6910w(0) <= x_prenodetwo_9_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6913w(0) <= x_prenodetwo_9_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6916w(0) <= x_prenodetwo_9_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6919w(0) <= x_prenodetwo_9_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6922w(0) <= x_prenodetwo_9_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6925w(0) <= x_prenodetwo_9_w(9);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7788w(0) <= y_prenode_10_w(0);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7869w(0) <= y_prenode_10_w(10);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7877w(0) <= y_prenode_10_w(11);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7885w(0) <= y_prenode_10_w(12);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7893w(0) <= y_prenode_10_w(13);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7901w(0) <= y_prenode_10_w(14);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7909w(0) <= y_prenode_10_w(15);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7917w(0) <= y_prenode_10_w(16);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7925w(0) <= y_prenode_10_w(17);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7933w(0) <= y_prenode_10_w(18);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7941w(0) <= y_prenode_10_w(19);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7797w(0) <= y_prenode_10_w(1);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7949w(0) <= y_prenode_10_w(20);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7957w(0) <= y_prenode_10_w(21);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7965w(0) <= y_prenode_10_w(22);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7973w(0) <= y_prenode_10_w(23);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7981w(0) <= y_prenode_10_w(24);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7989w(0) <= y_prenode_10_w(25);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7997w(0) <= y_prenode_10_w(26);
	wire_ccc_cordic_m_w_y_prenode_10_w_range8005w(0) <= y_prenode_10_w(27);
	wire_ccc_cordic_m_w_y_prenode_10_w_range8013w(0) <= y_prenode_10_w(28);
	wire_ccc_cordic_m_w_y_prenode_10_w_range8021w(0) <= y_prenode_10_w(29);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7805w(0) <= y_prenode_10_w(2);
	wire_ccc_cordic_m_w_y_prenode_10_w_range8029w(0) <= y_prenode_10_w(30);
	wire_ccc_cordic_m_w_y_prenode_10_w_range8037w(0) <= y_prenode_10_w(31);
	wire_ccc_cordic_m_w_y_prenode_10_w_range8045w(0) <= y_prenode_10_w(32);
	wire_ccc_cordic_m_w_y_prenode_10_w_range8053w(0) <= y_prenode_10_w(33);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7813w(0) <= y_prenode_10_w(3);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7821w(0) <= y_prenode_10_w(4);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7829w(0) <= y_prenode_10_w(5);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7837w(0) <= y_prenode_10_w(6);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7845w(0) <= y_prenode_10_w(7);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7853w(0) <= y_prenode_10_w(8);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7861w(0) <= y_prenode_10_w(9);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8595w(0) <= y_prenode_11_w(0);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8676w(0) <= y_prenode_11_w(10);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8684w(0) <= y_prenode_11_w(11);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8692w(0) <= y_prenode_11_w(12);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8700w(0) <= y_prenode_11_w(13);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8708w(0) <= y_prenode_11_w(14);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8716w(0) <= y_prenode_11_w(15);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8724w(0) <= y_prenode_11_w(16);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8732w(0) <= y_prenode_11_w(17);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8740w(0) <= y_prenode_11_w(18);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8748w(0) <= y_prenode_11_w(19);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8604w(0) <= y_prenode_11_w(1);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8756w(0) <= y_prenode_11_w(20);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8764w(0) <= y_prenode_11_w(21);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8772w(0) <= y_prenode_11_w(22);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8780w(0) <= y_prenode_11_w(23);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8788w(0) <= y_prenode_11_w(24);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8796w(0) <= y_prenode_11_w(25);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8804w(0) <= y_prenode_11_w(26);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8812w(0) <= y_prenode_11_w(27);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8820w(0) <= y_prenode_11_w(28);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8828w(0) <= y_prenode_11_w(29);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8612w(0) <= y_prenode_11_w(2);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8836w(0) <= y_prenode_11_w(30);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8844w(0) <= y_prenode_11_w(31);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8852w(0) <= y_prenode_11_w(32);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8860w(0) <= y_prenode_11_w(33);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8620w(0) <= y_prenode_11_w(3);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8628w(0) <= y_prenode_11_w(4);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8636w(0) <= y_prenode_11_w(5);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8644w(0) <= y_prenode_11_w(6);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8652w(0) <= y_prenode_11_w(7);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8660w(0) <= y_prenode_11_w(8);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8668w(0) <= y_prenode_11_w(9);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9397w(0) <= y_prenode_12_w(0);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9478w(0) <= y_prenode_12_w(10);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9486w(0) <= y_prenode_12_w(11);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9494w(0) <= y_prenode_12_w(12);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9502w(0) <= y_prenode_12_w(13);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9510w(0) <= y_prenode_12_w(14);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9518w(0) <= y_prenode_12_w(15);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9526w(0) <= y_prenode_12_w(16);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9534w(0) <= y_prenode_12_w(17);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9542w(0) <= y_prenode_12_w(18);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9550w(0) <= y_prenode_12_w(19);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9406w(0) <= y_prenode_12_w(1);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9558w(0) <= y_prenode_12_w(20);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9566w(0) <= y_prenode_12_w(21);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9574w(0) <= y_prenode_12_w(22);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9582w(0) <= y_prenode_12_w(23);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9590w(0) <= y_prenode_12_w(24);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9598w(0) <= y_prenode_12_w(25);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9606w(0) <= y_prenode_12_w(26);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9614w(0) <= y_prenode_12_w(27);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9622w(0) <= y_prenode_12_w(28);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9630w(0) <= y_prenode_12_w(29);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9414w(0) <= y_prenode_12_w(2);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9638w(0) <= y_prenode_12_w(30);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9646w(0) <= y_prenode_12_w(31);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9654w(0) <= y_prenode_12_w(32);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9662w(0) <= y_prenode_12_w(33);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9422w(0) <= y_prenode_12_w(3);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9430w(0) <= y_prenode_12_w(4);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9438w(0) <= y_prenode_12_w(5);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9446w(0) <= y_prenode_12_w(6);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9454w(0) <= y_prenode_12_w(7);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9462w(0) <= y_prenode_12_w(8);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9470w(0) <= y_prenode_12_w(9);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10194w(0) <= y_prenode_13_w(0);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10275w(0) <= y_prenode_13_w(10);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10283w(0) <= y_prenode_13_w(11);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10291w(0) <= y_prenode_13_w(12);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10299w(0) <= y_prenode_13_w(13);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10307w(0) <= y_prenode_13_w(14);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10315w(0) <= y_prenode_13_w(15);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10323w(0) <= y_prenode_13_w(16);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10331w(0) <= y_prenode_13_w(17);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10339w(0) <= y_prenode_13_w(18);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10347w(0) <= y_prenode_13_w(19);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10203w(0) <= y_prenode_13_w(1);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10355w(0) <= y_prenode_13_w(20);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10363w(0) <= y_prenode_13_w(21);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10371w(0) <= y_prenode_13_w(22);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10379w(0) <= y_prenode_13_w(23);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10387w(0) <= y_prenode_13_w(24);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10395w(0) <= y_prenode_13_w(25);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10403w(0) <= y_prenode_13_w(26);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10411w(0) <= y_prenode_13_w(27);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10419w(0) <= y_prenode_13_w(28);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10427w(0) <= y_prenode_13_w(29);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10211w(0) <= y_prenode_13_w(2);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10435w(0) <= y_prenode_13_w(30);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10443w(0) <= y_prenode_13_w(31);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10451w(0) <= y_prenode_13_w(32);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10459w(0) <= y_prenode_13_w(33);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10219w(0) <= y_prenode_13_w(3);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10227w(0) <= y_prenode_13_w(4);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10235w(0) <= y_prenode_13_w(5);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10243w(0) <= y_prenode_13_w(6);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10251w(0) <= y_prenode_13_w(7);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10259w(0) <= y_prenode_13_w(8);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10267w(0) <= y_prenode_13_w(9);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1152w(0) <= y_prenode_2_w(0);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1233w(0) <= y_prenode_2_w(10);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1241w(0) <= y_prenode_2_w(11);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1249w(0) <= y_prenode_2_w(12);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1257w(0) <= y_prenode_2_w(13);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1265w(0) <= y_prenode_2_w(14);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1273w(0) <= y_prenode_2_w(15);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1281w(0) <= y_prenode_2_w(16);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1289w(0) <= y_prenode_2_w(17);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1297w(0) <= y_prenode_2_w(18);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1305w(0) <= y_prenode_2_w(19);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1161w(0) <= y_prenode_2_w(1);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1313w(0) <= y_prenode_2_w(20);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1321w(0) <= y_prenode_2_w(21);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1329w(0) <= y_prenode_2_w(22);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1337w(0) <= y_prenode_2_w(23);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1345w(0) <= y_prenode_2_w(24);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1353w(0) <= y_prenode_2_w(25);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1361w(0) <= y_prenode_2_w(26);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1369w(0) <= y_prenode_2_w(27);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1377w(0) <= y_prenode_2_w(28);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1385w(0) <= y_prenode_2_w(29);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1169w(0) <= y_prenode_2_w(2);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1393w(0) <= y_prenode_2_w(30);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1401w(0) <= y_prenode_2_w(31);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1409w(0) <= y_prenode_2_w(32);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1417w(0) <= y_prenode_2_w(33);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1177w(0) <= y_prenode_2_w(3);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1185w(0) <= y_prenode_2_w(4);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1193w(0) <= y_prenode_2_w(5);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1201w(0) <= y_prenode_2_w(6);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1209w(0) <= y_prenode_2_w(7);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1217w(0) <= y_prenode_2_w(8);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1225w(0) <= y_prenode_2_w(9);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1999w(0) <= y_prenode_3_w(0);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2080w(0) <= y_prenode_3_w(10);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2088w(0) <= y_prenode_3_w(11);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2096w(0) <= y_prenode_3_w(12);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2104w(0) <= y_prenode_3_w(13);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2112w(0) <= y_prenode_3_w(14);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2120w(0) <= y_prenode_3_w(15);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2128w(0) <= y_prenode_3_w(16);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2136w(0) <= y_prenode_3_w(17);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2144w(0) <= y_prenode_3_w(18);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2152w(0) <= y_prenode_3_w(19);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2008w(0) <= y_prenode_3_w(1);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2160w(0) <= y_prenode_3_w(20);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2168w(0) <= y_prenode_3_w(21);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2176w(0) <= y_prenode_3_w(22);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2184w(0) <= y_prenode_3_w(23);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2192w(0) <= y_prenode_3_w(24);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2200w(0) <= y_prenode_3_w(25);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2208w(0) <= y_prenode_3_w(26);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2216w(0) <= y_prenode_3_w(27);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2224w(0) <= y_prenode_3_w(28);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2232w(0) <= y_prenode_3_w(29);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2016w(0) <= y_prenode_3_w(2);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2240w(0) <= y_prenode_3_w(30);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2248w(0) <= y_prenode_3_w(31);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2256w(0) <= y_prenode_3_w(32);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2264w(0) <= y_prenode_3_w(33);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2024w(0) <= y_prenode_3_w(3);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2032w(0) <= y_prenode_3_w(4);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2040w(0) <= y_prenode_3_w(5);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2048w(0) <= y_prenode_3_w(6);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2056w(0) <= y_prenode_3_w(7);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2064w(0) <= y_prenode_3_w(8);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2072w(0) <= y_prenode_3_w(9);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2841w(0) <= y_prenode_4_w(0);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2922w(0) <= y_prenode_4_w(10);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2930w(0) <= y_prenode_4_w(11);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2938w(0) <= y_prenode_4_w(12);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2946w(0) <= y_prenode_4_w(13);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2954w(0) <= y_prenode_4_w(14);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2962w(0) <= y_prenode_4_w(15);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2970w(0) <= y_prenode_4_w(16);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2978w(0) <= y_prenode_4_w(17);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2986w(0) <= y_prenode_4_w(18);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2994w(0) <= y_prenode_4_w(19);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2850w(0) <= y_prenode_4_w(1);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3002w(0) <= y_prenode_4_w(20);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3010w(0) <= y_prenode_4_w(21);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3018w(0) <= y_prenode_4_w(22);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3026w(0) <= y_prenode_4_w(23);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3034w(0) <= y_prenode_4_w(24);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3042w(0) <= y_prenode_4_w(25);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3050w(0) <= y_prenode_4_w(26);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3058w(0) <= y_prenode_4_w(27);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3066w(0) <= y_prenode_4_w(28);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3074w(0) <= y_prenode_4_w(29);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2858w(0) <= y_prenode_4_w(2);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3082w(0) <= y_prenode_4_w(30);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3090w(0) <= y_prenode_4_w(31);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3098w(0) <= y_prenode_4_w(32);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3106w(0) <= y_prenode_4_w(33);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2866w(0) <= y_prenode_4_w(3);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2874w(0) <= y_prenode_4_w(4);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2882w(0) <= y_prenode_4_w(5);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2890w(0) <= y_prenode_4_w(6);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2898w(0) <= y_prenode_4_w(7);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2906w(0) <= y_prenode_4_w(8);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2914w(0) <= y_prenode_4_w(9);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3678w(0) <= y_prenode_5_w(0);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3759w(0) <= y_prenode_5_w(10);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3767w(0) <= y_prenode_5_w(11);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3775w(0) <= y_prenode_5_w(12);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3783w(0) <= y_prenode_5_w(13);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3791w(0) <= y_prenode_5_w(14);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3799w(0) <= y_prenode_5_w(15);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3807w(0) <= y_prenode_5_w(16);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3815w(0) <= y_prenode_5_w(17);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3823w(0) <= y_prenode_5_w(18);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3831w(0) <= y_prenode_5_w(19);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3687w(0) <= y_prenode_5_w(1);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3839w(0) <= y_prenode_5_w(20);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3847w(0) <= y_prenode_5_w(21);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3855w(0) <= y_prenode_5_w(22);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3863w(0) <= y_prenode_5_w(23);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3871w(0) <= y_prenode_5_w(24);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3879w(0) <= y_prenode_5_w(25);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3887w(0) <= y_prenode_5_w(26);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3895w(0) <= y_prenode_5_w(27);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3903w(0) <= y_prenode_5_w(28);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3911w(0) <= y_prenode_5_w(29);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3695w(0) <= y_prenode_5_w(2);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3919w(0) <= y_prenode_5_w(30);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3927w(0) <= y_prenode_5_w(31);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3935w(0) <= y_prenode_5_w(32);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3943w(0) <= y_prenode_5_w(33);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3703w(0) <= y_prenode_5_w(3);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3711w(0) <= y_prenode_5_w(4);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3719w(0) <= y_prenode_5_w(5);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3727w(0) <= y_prenode_5_w(6);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3735w(0) <= y_prenode_5_w(7);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3743w(0) <= y_prenode_5_w(8);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3751w(0) <= y_prenode_5_w(9);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4510w(0) <= y_prenode_6_w(0);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4591w(0) <= y_prenode_6_w(10);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4599w(0) <= y_prenode_6_w(11);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4607w(0) <= y_prenode_6_w(12);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4615w(0) <= y_prenode_6_w(13);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4623w(0) <= y_prenode_6_w(14);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4631w(0) <= y_prenode_6_w(15);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4639w(0) <= y_prenode_6_w(16);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4647w(0) <= y_prenode_6_w(17);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4655w(0) <= y_prenode_6_w(18);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4663w(0) <= y_prenode_6_w(19);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4519w(0) <= y_prenode_6_w(1);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4671w(0) <= y_prenode_6_w(20);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4679w(0) <= y_prenode_6_w(21);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4687w(0) <= y_prenode_6_w(22);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4695w(0) <= y_prenode_6_w(23);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4703w(0) <= y_prenode_6_w(24);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4711w(0) <= y_prenode_6_w(25);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4719w(0) <= y_prenode_6_w(26);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4727w(0) <= y_prenode_6_w(27);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4735w(0) <= y_prenode_6_w(28);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4743w(0) <= y_prenode_6_w(29);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4527w(0) <= y_prenode_6_w(2);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4751w(0) <= y_prenode_6_w(30);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4759w(0) <= y_prenode_6_w(31);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4767w(0) <= y_prenode_6_w(32);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4775w(0) <= y_prenode_6_w(33);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4535w(0) <= y_prenode_6_w(3);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4543w(0) <= y_prenode_6_w(4);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4551w(0) <= y_prenode_6_w(5);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4559w(0) <= y_prenode_6_w(6);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4567w(0) <= y_prenode_6_w(7);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4575w(0) <= y_prenode_6_w(8);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4583w(0) <= y_prenode_6_w(9);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5337w(0) <= y_prenode_7_w(0);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5418w(0) <= y_prenode_7_w(10);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5426w(0) <= y_prenode_7_w(11);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5434w(0) <= y_prenode_7_w(12);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5442w(0) <= y_prenode_7_w(13);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5450w(0) <= y_prenode_7_w(14);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5458w(0) <= y_prenode_7_w(15);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5466w(0) <= y_prenode_7_w(16);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5474w(0) <= y_prenode_7_w(17);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5482w(0) <= y_prenode_7_w(18);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5490w(0) <= y_prenode_7_w(19);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5346w(0) <= y_prenode_7_w(1);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5498w(0) <= y_prenode_7_w(20);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5506w(0) <= y_prenode_7_w(21);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5514w(0) <= y_prenode_7_w(22);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5522w(0) <= y_prenode_7_w(23);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5530w(0) <= y_prenode_7_w(24);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5538w(0) <= y_prenode_7_w(25);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5546w(0) <= y_prenode_7_w(26);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5554w(0) <= y_prenode_7_w(27);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5562w(0) <= y_prenode_7_w(28);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5570w(0) <= y_prenode_7_w(29);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5354w(0) <= y_prenode_7_w(2);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5578w(0) <= y_prenode_7_w(30);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5586w(0) <= y_prenode_7_w(31);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5594w(0) <= y_prenode_7_w(32);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5602w(0) <= y_prenode_7_w(33);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5362w(0) <= y_prenode_7_w(3);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5370w(0) <= y_prenode_7_w(4);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5378w(0) <= y_prenode_7_w(5);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5386w(0) <= y_prenode_7_w(6);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5394w(0) <= y_prenode_7_w(7);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5402w(0) <= y_prenode_7_w(8);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5410w(0) <= y_prenode_7_w(9);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6159w(0) <= y_prenode_8_w(0);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6240w(0) <= y_prenode_8_w(10);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6248w(0) <= y_prenode_8_w(11);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6256w(0) <= y_prenode_8_w(12);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6264w(0) <= y_prenode_8_w(13);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6272w(0) <= y_prenode_8_w(14);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6280w(0) <= y_prenode_8_w(15);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6288w(0) <= y_prenode_8_w(16);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6296w(0) <= y_prenode_8_w(17);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6304w(0) <= y_prenode_8_w(18);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6312w(0) <= y_prenode_8_w(19);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6168w(0) <= y_prenode_8_w(1);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6320w(0) <= y_prenode_8_w(20);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6328w(0) <= y_prenode_8_w(21);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6336w(0) <= y_prenode_8_w(22);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6344w(0) <= y_prenode_8_w(23);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6352w(0) <= y_prenode_8_w(24);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6360w(0) <= y_prenode_8_w(25);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6368w(0) <= y_prenode_8_w(26);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6376w(0) <= y_prenode_8_w(27);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6384w(0) <= y_prenode_8_w(28);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6392w(0) <= y_prenode_8_w(29);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6176w(0) <= y_prenode_8_w(2);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6400w(0) <= y_prenode_8_w(30);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6408w(0) <= y_prenode_8_w(31);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6416w(0) <= y_prenode_8_w(32);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6424w(0) <= y_prenode_8_w(33);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6184w(0) <= y_prenode_8_w(3);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6192w(0) <= y_prenode_8_w(4);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6200w(0) <= y_prenode_8_w(5);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6208w(0) <= y_prenode_8_w(6);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6216w(0) <= y_prenode_8_w(7);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6224w(0) <= y_prenode_8_w(8);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6232w(0) <= y_prenode_8_w(9);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6976w(0) <= y_prenode_9_w(0);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7057w(0) <= y_prenode_9_w(10);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7065w(0) <= y_prenode_9_w(11);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7073w(0) <= y_prenode_9_w(12);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7081w(0) <= y_prenode_9_w(13);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7089w(0) <= y_prenode_9_w(14);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7097w(0) <= y_prenode_9_w(15);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7105w(0) <= y_prenode_9_w(16);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7113w(0) <= y_prenode_9_w(17);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7121w(0) <= y_prenode_9_w(18);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7129w(0) <= y_prenode_9_w(19);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6985w(0) <= y_prenode_9_w(1);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7137w(0) <= y_prenode_9_w(20);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7145w(0) <= y_prenode_9_w(21);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7153w(0) <= y_prenode_9_w(22);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7161w(0) <= y_prenode_9_w(23);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7169w(0) <= y_prenode_9_w(24);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7177w(0) <= y_prenode_9_w(25);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7185w(0) <= y_prenode_9_w(26);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7193w(0) <= y_prenode_9_w(27);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7201w(0) <= y_prenode_9_w(28);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7209w(0) <= y_prenode_9_w(29);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6993w(0) <= y_prenode_9_w(2);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7217w(0) <= y_prenode_9_w(30);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7225w(0) <= y_prenode_9_w(31);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7233w(0) <= y_prenode_9_w(32);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7241w(0) <= y_prenode_9_w(33);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7001w(0) <= y_prenode_9_w(3);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7009w(0) <= y_prenode_9_w(4);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7017w(0) <= y_prenode_9_w(5);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7025w(0) <= y_prenode_9_w(6);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7033w(0) <= y_prenode_9_w(7);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7041w(0) <= y_prenode_9_w(8);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7049w(0) <= y_prenode_9_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7572w(0) <= y_prenodeone_10_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7631w(0) <= y_prenodeone_10_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7637w(0) <= y_prenodeone_10_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7643w(0) <= y_prenodeone_10_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7649w(0) <= y_prenodeone_10_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7655w(0) <= y_prenodeone_10_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7661w(0) <= y_prenodeone_10_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7667w(0) <= y_prenodeone_10_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7673w(0) <= y_prenodeone_10_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7679w(0) <= y_prenodeone_10_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7685w(0) <= y_prenodeone_10_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7577w(0) <= y_prenodeone_10_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7691w(0) <= y_prenodeone_10_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7697w(0) <= y_prenodeone_10_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7703w(0) <= y_prenodeone_10_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7709w(0) <= y_prenodeone_10_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7712w(0) <= y_prenodeone_10_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7526w(0) <= y_prenodeone_10_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7529w(0) <= y_prenodeone_10_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7531w(0) <= y_prenodeone_10_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7533w(0) <= y_prenodeone_10_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7535w(0) <= y_prenodeone_10_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7583w(0) <= y_prenodeone_10_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7537w(0) <= y_prenodeone_10_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7539w(0) <= y_prenodeone_10_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7541w(0) <= y_prenodeone_10_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7543w(0) <= y_prenodeone_10_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7589w(0) <= y_prenodeone_10_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7595w(0) <= y_prenodeone_10_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7601w(0) <= y_prenodeone_10_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7607w(0) <= y_prenodeone_10_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7613w(0) <= y_prenodeone_10_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7619w(0) <= y_prenodeone_10_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7625w(0) <= y_prenodeone_10_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8388w(0) <= y_prenodeone_11_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8447w(0) <= y_prenodeone_11_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8453w(0) <= y_prenodeone_11_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8459w(0) <= y_prenodeone_11_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8465w(0) <= y_prenodeone_11_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8471w(0) <= y_prenodeone_11_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8477w(0) <= y_prenodeone_11_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8483w(0) <= y_prenodeone_11_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8489w(0) <= y_prenodeone_11_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8495w(0) <= y_prenodeone_11_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8501w(0) <= y_prenodeone_11_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8393w(0) <= y_prenodeone_11_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8507w(0) <= y_prenodeone_11_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8513w(0) <= y_prenodeone_11_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8519w(0) <= y_prenodeone_11_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8522w(0) <= y_prenodeone_11_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8338w(0) <= y_prenodeone_11_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8341w(0) <= y_prenodeone_11_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8343w(0) <= y_prenodeone_11_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8345w(0) <= y_prenodeone_11_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8347w(0) <= y_prenodeone_11_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8349w(0) <= y_prenodeone_11_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8399w(0) <= y_prenodeone_11_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8351w(0) <= y_prenodeone_11_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8353w(0) <= y_prenodeone_11_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8355w(0) <= y_prenodeone_11_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8357w(0) <= y_prenodeone_11_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8405w(0) <= y_prenodeone_11_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8411w(0) <= y_prenodeone_11_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8417w(0) <= y_prenodeone_11_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8423w(0) <= y_prenodeone_11_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8429w(0) <= y_prenodeone_11_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8435w(0) <= y_prenodeone_11_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8441w(0) <= y_prenodeone_11_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9199w(0) <= y_prenodeone_12_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9258w(0) <= y_prenodeone_12_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9264w(0) <= y_prenodeone_12_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9270w(0) <= y_prenodeone_12_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9276w(0) <= y_prenodeone_12_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9282w(0) <= y_prenodeone_12_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9288w(0) <= y_prenodeone_12_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9294w(0) <= y_prenodeone_12_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9300w(0) <= y_prenodeone_12_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9306w(0) <= y_prenodeone_12_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9312w(0) <= y_prenodeone_12_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9204w(0) <= y_prenodeone_12_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9318w(0) <= y_prenodeone_12_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9324w(0) <= y_prenodeone_12_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9327w(0) <= y_prenodeone_12_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9145w(0) <= y_prenodeone_12_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9148w(0) <= y_prenodeone_12_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9150w(0) <= y_prenodeone_12_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9152w(0) <= y_prenodeone_12_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9154w(0) <= y_prenodeone_12_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9156w(0) <= y_prenodeone_12_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9158w(0) <= y_prenodeone_12_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9210w(0) <= y_prenodeone_12_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9160w(0) <= y_prenodeone_12_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9162w(0) <= y_prenodeone_12_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9164w(0) <= y_prenodeone_12_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9166w(0) <= y_prenodeone_12_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9216w(0) <= y_prenodeone_12_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9222w(0) <= y_prenodeone_12_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9228w(0) <= y_prenodeone_12_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9234w(0) <= y_prenodeone_12_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9240w(0) <= y_prenodeone_12_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9246w(0) <= y_prenodeone_12_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9252w(0) <= y_prenodeone_12_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10005w(0) <= y_prenodeone_13_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10064w(0) <= y_prenodeone_13_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10070w(0) <= y_prenodeone_13_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10076w(0) <= y_prenodeone_13_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10082w(0) <= y_prenodeone_13_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10088w(0) <= y_prenodeone_13_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10094w(0) <= y_prenodeone_13_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10100w(0) <= y_prenodeone_13_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10106w(0) <= y_prenodeone_13_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10112w(0) <= y_prenodeone_13_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10118w(0) <= y_prenodeone_13_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10010w(0) <= y_prenodeone_13_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10124w(0) <= y_prenodeone_13_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10127w(0) <= y_prenodeone_13_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9947w(0) <= y_prenodeone_13_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9950w(0) <= y_prenodeone_13_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9952w(0) <= y_prenodeone_13_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9954w(0) <= y_prenodeone_13_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9956w(0) <= y_prenodeone_13_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9958w(0) <= y_prenodeone_13_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9960w(0) <= y_prenodeone_13_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9962w(0) <= y_prenodeone_13_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10016w(0) <= y_prenodeone_13_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9964w(0) <= y_prenodeone_13_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9966w(0) <= y_prenodeone_13_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9968w(0) <= y_prenodeone_13_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9970w(0) <= y_prenodeone_13_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10022w(0) <= y_prenodeone_13_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10028w(0) <= y_prenodeone_13_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10034w(0) <= y_prenodeone_13_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10040w(0) <= y_prenodeone_13_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10046w(0) <= y_prenodeone_13_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10052w(0) <= y_prenodeone_13_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10058w(0) <= y_prenodeone_13_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range864w(0) <= y_prenodeone_2_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range923w(0) <= y_prenodeone_2_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range929w(0) <= y_prenodeone_2_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range935w(0) <= y_prenodeone_2_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range941w(0) <= y_prenodeone_2_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range947w(0) <= y_prenodeone_2_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range953w(0) <= y_prenodeone_2_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range959w(0) <= y_prenodeone_2_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range965w(0) <= y_prenodeone_2_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range971w(0) <= y_prenodeone_2_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range977w(0) <= y_prenodeone_2_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range869w(0) <= y_prenodeone_2_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range983w(0) <= y_prenodeone_2_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range989w(0) <= y_prenodeone_2_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range995w(0) <= y_prenodeone_2_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range1001w(0) <= y_prenodeone_2_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range1007w(0) <= y_prenodeone_2_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range1013w(0) <= y_prenodeone_2_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range1019w(0) <= y_prenodeone_2_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range1025w(0) <= y_prenodeone_2_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range1031w(0) <= y_prenodeone_2_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range1037w(0) <= y_prenodeone_2_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range875w(0) <= y_prenodeone_2_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range1043w(0) <= y_prenodeone_2_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range1049w(0) <= y_prenodeone_2_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range1052w(0) <= y_prenodeone_2_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range850w(0) <= y_prenodeone_2_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range881w(0) <= y_prenodeone_2_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range887w(0) <= y_prenodeone_2_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range893w(0) <= y_prenodeone_2_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range899w(0) <= y_prenodeone_2_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range905w(0) <= y_prenodeone_2_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range911w(0) <= y_prenodeone_2_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range917w(0) <= y_prenodeone_2_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1720w(0) <= y_prenodeone_3_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1779w(0) <= y_prenodeone_3_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1785w(0) <= y_prenodeone_3_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1791w(0) <= y_prenodeone_3_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1797w(0) <= y_prenodeone_3_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1803w(0) <= y_prenodeone_3_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1809w(0) <= y_prenodeone_3_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1815w(0) <= y_prenodeone_3_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1821w(0) <= y_prenodeone_3_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1827w(0) <= y_prenodeone_3_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1833w(0) <= y_prenodeone_3_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1725w(0) <= y_prenodeone_3_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1839w(0) <= y_prenodeone_3_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1845w(0) <= y_prenodeone_3_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1851w(0) <= y_prenodeone_3_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1857w(0) <= y_prenodeone_3_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1863w(0) <= y_prenodeone_3_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1869w(0) <= y_prenodeone_3_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1875w(0) <= y_prenodeone_3_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1881w(0) <= y_prenodeone_3_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1887w(0) <= y_prenodeone_3_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1893w(0) <= y_prenodeone_3_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1731w(0) <= y_prenodeone_3_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1899w(0) <= y_prenodeone_3_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1902w(0) <= y_prenodeone_3_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1702w(0) <= y_prenodeone_3_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1705w(0) <= y_prenodeone_3_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1737w(0) <= y_prenodeone_3_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1743w(0) <= y_prenodeone_3_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1749w(0) <= y_prenodeone_3_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1755w(0) <= y_prenodeone_3_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1761w(0) <= y_prenodeone_3_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1767w(0) <= y_prenodeone_3_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1773w(0) <= y_prenodeone_3_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2571w(0) <= y_prenodeone_4_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2630w(0) <= y_prenodeone_4_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2636w(0) <= y_prenodeone_4_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2642w(0) <= y_prenodeone_4_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2648w(0) <= y_prenodeone_4_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2654w(0) <= y_prenodeone_4_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2660w(0) <= y_prenodeone_4_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2666w(0) <= y_prenodeone_4_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2672w(0) <= y_prenodeone_4_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2678w(0) <= y_prenodeone_4_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2684w(0) <= y_prenodeone_4_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2576w(0) <= y_prenodeone_4_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2690w(0) <= y_prenodeone_4_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2696w(0) <= y_prenodeone_4_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2702w(0) <= y_prenodeone_4_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2708w(0) <= y_prenodeone_4_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2714w(0) <= y_prenodeone_4_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2720w(0) <= y_prenodeone_4_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2726w(0) <= y_prenodeone_4_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2732w(0) <= y_prenodeone_4_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2738w(0) <= y_prenodeone_4_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2744w(0) <= y_prenodeone_4_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2582w(0) <= y_prenodeone_4_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2747w(0) <= y_prenodeone_4_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2549w(0) <= y_prenodeone_4_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2552w(0) <= y_prenodeone_4_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2554w(0) <= y_prenodeone_4_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2588w(0) <= y_prenodeone_4_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2594w(0) <= y_prenodeone_4_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2600w(0) <= y_prenodeone_4_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2606w(0) <= y_prenodeone_4_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2612w(0) <= y_prenodeone_4_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2618w(0) <= y_prenodeone_4_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2624w(0) <= y_prenodeone_4_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3417w(0) <= y_prenodeone_5_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3476w(0) <= y_prenodeone_5_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3482w(0) <= y_prenodeone_5_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3488w(0) <= y_prenodeone_5_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3494w(0) <= y_prenodeone_5_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3500w(0) <= y_prenodeone_5_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3506w(0) <= y_prenodeone_5_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3512w(0) <= y_prenodeone_5_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3518w(0) <= y_prenodeone_5_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3524w(0) <= y_prenodeone_5_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3530w(0) <= y_prenodeone_5_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3422w(0) <= y_prenodeone_5_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3536w(0) <= y_prenodeone_5_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3542w(0) <= y_prenodeone_5_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3548w(0) <= y_prenodeone_5_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3554w(0) <= y_prenodeone_5_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3560w(0) <= y_prenodeone_5_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3566w(0) <= y_prenodeone_5_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3572w(0) <= y_prenodeone_5_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3578w(0) <= y_prenodeone_5_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3584w(0) <= y_prenodeone_5_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3587w(0) <= y_prenodeone_5_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3428w(0) <= y_prenodeone_5_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3391w(0) <= y_prenodeone_5_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3394w(0) <= y_prenodeone_5_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3396w(0) <= y_prenodeone_5_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3398w(0) <= y_prenodeone_5_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3434w(0) <= y_prenodeone_5_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3440w(0) <= y_prenodeone_5_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3446w(0) <= y_prenodeone_5_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3452w(0) <= y_prenodeone_5_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3458w(0) <= y_prenodeone_5_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3464w(0) <= y_prenodeone_5_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3470w(0) <= y_prenodeone_5_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4258w(0) <= y_prenodeone_6_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4317w(0) <= y_prenodeone_6_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4323w(0) <= y_prenodeone_6_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4329w(0) <= y_prenodeone_6_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4335w(0) <= y_prenodeone_6_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4341w(0) <= y_prenodeone_6_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4347w(0) <= y_prenodeone_6_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4353w(0) <= y_prenodeone_6_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4359w(0) <= y_prenodeone_6_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4365w(0) <= y_prenodeone_6_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4371w(0) <= y_prenodeone_6_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4263w(0) <= y_prenodeone_6_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4377w(0) <= y_prenodeone_6_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4383w(0) <= y_prenodeone_6_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4389w(0) <= y_prenodeone_6_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4395w(0) <= y_prenodeone_6_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4401w(0) <= y_prenodeone_6_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4407w(0) <= y_prenodeone_6_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4413w(0) <= y_prenodeone_6_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4419w(0) <= y_prenodeone_6_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4422w(0) <= y_prenodeone_6_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4228w(0) <= y_prenodeone_6_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4269w(0) <= y_prenodeone_6_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4231w(0) <= y_prenodeone_6_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4233w(0) <= y_prenodeone_6_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4235w(0) <= y_prenodeone_6_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4237w(0) <= y_prenodeone_6_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4275w(0) <= y_prenodeone_6_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4281w(0) <= y_prenodeone_6_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4287w(0) <= y_prenodeone_6_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4293w(0) <= y_prenodeone_6_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4299w(0) <= y_prenodeone_6_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4305w(0) <= y_prenodeone_6_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4311w(0) <= y_prenodeone_6_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5094w(0) <= y_prenodeone_7_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5153w(0) <= y_prenodeone_7_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5159w(0) <= y_prenodeone_7_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5165w(0) <= y_prenodeone_7_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5171w(0) <= y_prenodeone_7_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5177w(0) <= y_prenodeone_7_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5183w(0) <= y_prenodeone_7_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5189w(0) <= y_prenodeone_7_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5195w(0) <= y_prenodeone_7_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5201w(0) <= y_prenodeone_7_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5207w(0) <= y_prenodeone_7_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5099w(0) <= y_prenodeone_7_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5213w(0) <= y_prenodeone_7_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5219w(0) <= y_prenodeone_7_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5225w(0) <= y_prenodeone_7_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5231w(0) <= y_prenodeone_7_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5237w(0) <= y_prenodeone_7_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5243w(0) <= y_prenodeone_7_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5249w(0) <= y_prenodeone_7_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5252w(0) <= y_prenodeone_7_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5060w(0) <= y_prenodeone_7_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5063w(0) <= y_prenodeone_7_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5105w(0) <= y_prenodeone_7_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5065w(0) <= y_prenodeone_7_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5067w(0) <= y_prenodeone_7_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5069w(0) <= y_prenodeone_7_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5071w(0) <= y_prenodeone_7_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5111w(0) <= y_prenodeone_7_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5117w(0) <= y_prenodeone_7_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5123w(0) <= y_prenodeone_7_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5129w(0) <= y_prenodeone_7_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5135w(0) <= y_prenodeone_7_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5141w(0) <= y_prenodeone_7_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5147w(0) <= y_prenodeone_7_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5925w(0) <= y_prenodeone_8_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5984w(0) <= y_prenodeone_8_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5990w(0) <= y_prenodeone_8_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5996w(0) <= y_prenodeone_8_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6002w(0) <= y_prenodeone_8_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6008w(0) <= y_prenodeone_8_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6014w(0) <= y_prenodeone_8_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6020w(0) <= y_prenodeone_8_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6026w(0) <= y_prenodeone_8_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6032w(0) <= y_prenodeone_8_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6038w(0) <= y_prenodeone_8_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5930w(0) <= y_prenodeone_8_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6044w(0) <= y_prenodeone_8_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6050w(0) <= y_prenodeone_8_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6056w(0) <= y_prenodeone_8_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6062w(0) <= y_prenodeone_8_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6068w(0) <= y_prenodeone_8_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6074w(0) <= y_prenodeone_8_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6077w(0) <= y_prenodeone_8_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5887w(0) <= y_prenodeone_8_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5890w(0) <= y_prenodeone_8_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5892w(0) <= y_prenodeone_8_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5936w(0) <= y_prenodeone_8_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5894w(0) <= y_prenodeone_8_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5896w(0) <= y_prenodeone_8_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5898w(0) <= y_prenodeone_8_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5900w(0) <= y_prenodeone_8_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5942w(0) <= y_prenodeone_8_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5948w(0) <= y_prenodeone_8_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5954w(0) <= y_prenodeone_8_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5960w(0) <= y_prenodeone_8_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5966w(0) <= y_prenodeone_8_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5972w(0) <= y_prenodeone_8_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5978w(0) <= y_prenodeone_8_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6751w(0) <= y_prenodeone_9_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6810w(0) <= y_prenodeone_9_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6816w(0) <= y_prenodeone_9_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6822w(0) <= y_prenodeone_9_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6828w(0) <= y_prenodeone_9_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6834w(0) <= y_prenodeone_9_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6840w(0) <= y_prenodeone_9_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6846w(0) <= y_prenodeone_9_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6852w(0) <= y_prenodeone_9_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6858w(0) <= y_prenodeone_9_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6864w(0) <= y_prenodeone_9_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6756w(0) <= y_prenodeone_9_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6870w(0) <= y_prenodeone_9_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6876w(0) <= y_prenodeone_9_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6882w(0) <= y_prenodeone_9_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6888w(0) <= y_prenodeone_9_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6894w(0) <= y_prenodeone_9_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6897w(0) <= y_prenodeone_9_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6709w(0) <= y_prenodeone_9_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6712w(0) <= y_prenodeone_9_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6714w(0) <= y_prenodeone_9_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6716w(0) <= y_prenodeone_9_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6762w(0) <= y_prenodeone_9_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6718w(0) <= y_prenodeone_9_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6720w(0) <= y_prenodeone_9_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6722w(0) <= y_prenodeone_9_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6724w(0) <= y_prenodeone_9_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6768w(0) <= y_prenodeone_9_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6774w(0) <= y_prenodeone_9_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6780w(0) <= y_prenodeone_9_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6786w(0) <= y_prenodeone_9_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6792w(0) <= y_prenodeone_9_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6798w(0) <= y_prenodeone_9_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6804w(0) <= y_prenodeone_9_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7715w(0) <= y_prenodetwo_10_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7744w(0) <= y_prenodetwo_10_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7747w(0) <= y_prenodetwo_10_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7750w(0) <= y_prenodetwo_10_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7753w(0) <= y_prenodetwo_10_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7756w(0) <= y_prenodetwo_10_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7759w(0) <= y_prenodetwo_10_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7762w(0) <= y_prenodetwo_10_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7765w(0) <= y_prenodetwo_10_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7768w(0) <= y_prenodetwo_10_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7771w(0) <= y_prenodetwo_10_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7717w(0) <= y_prenodetwo_10_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7774w(0) <= y_prenodetwo_10_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7777w(0) <= y_prenodetwo_10_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7780w(0) <= y_prenodetwo_10_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7546w(0) <= y_prenodetwo_10_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7549w(0) <= y_prenodetwo_10_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7551w(0) <= y_prenodetwo_10_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7553w(0) <= y_prenodetwo_10_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7555w(0) <= y_prenodetwo_10_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7557w(0) <= y_prenodetwo_10_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7559w(0) <= y_prenodetwo_10_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7720w(0) <= y_prenodetwo_10_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7561w(0) <= y_prenodetwo_10_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7563w(0) <= y_prenodetwo_10_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7565w(0) <= y_prenodetwo_10_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7567w(0) <= y_prenodetwo_10_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7723w(0) <= y_prenodetwo_10_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7726w(0) <= y_prenodetwo_10_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7729w(0) <= y_prenodetwo_10_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7732w(0) <= y_prenodetwo_10_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7735w(0) <= y_prenodetwo_10_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7738w(0) <= y_prenodetwo_10_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7741w(0) <= y_prenodetwo_10_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8525w(0) <= y_prenodetwo_11_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8554w(0) <= y_prenodetwo_11_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8557w(0) <= y_prenodetwo_11_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8560w(0) <= y_prenodetwo_11_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8563w(0) <= y_prenodetwo_11_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8566w(0) <= y_prenodetwo_11_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8569w(0) <= y_prenodetwo_11_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8572w(0) <= y_prenodetwo_11_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8575w(0) <= y_prenodetwo_11_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8578w(0) <= y_prenodetwo_11_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8581w(0) <= y_prenodetwo_11_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8527w(0) <= y_prenodetwo_11_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8584w(0) <= y_prenodetwo_11_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8587w(0) <= y_prenodetwo_11_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8360w(0) <= y_prenodetwo_11_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8363w(0) <= y_prenodetwo_11_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8365w(0) <= y_prenodetwo_11_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8367w(0) <= y_prenodetwo_11_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8369w(0) <= y_prenodetwo_11_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8371w(0) <= y_prenodetwo_11_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8373w(0) <= y_prenodetwo_11_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8375w(0) <= y_prenodetwo_11_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8530w(0) <= y_prenodetwo_11_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8377w(0) <= y_prenodetwo_11_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8379w(0) <= y_prenodetwo_11_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8381w(0) <= y_prenodetwo_11_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8383w(0) <= y_prenodetwo_11_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8533w(0) <= y_prenodetwo_11_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8536w(0) <= y_prenodetwo_11_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8539w(0) <= y_prenodetwo_11_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8542w(0) <= y_prenodetwo_11_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8545w(0) <= y_prenodetwo_11_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8548w(0) <= y_prenodetwo_11_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8551w(0) <= y_prenodetwo_11_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9330w(0) <= y_prenodetwo_12_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9359w(0) <= y_prenodetwo_12_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9362w(0) <= y_prenodetwo_12_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9365w(0) <= y_prenodetwo_12_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9368w(0) <= y_prenodetwo_12_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9371w(0) <= y_prenodetwo_12_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9374w(0) <= y_prenodetwo_12_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9377w(0) <= y_prenodetwo_12_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9380w(0) <= y_prenodetwo_12_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9383w(0) <= y_prenodetwo_12_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9386w(0) <= y_prenodetwo_12_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9332w(0) <= y_prenodetwo_12_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9389w(0) <= y_prenodetwo_12_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9169w(0) <= y_prenodetwo_12_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9172w(0) <= y_prenodetwo_12_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9174w(0) <= y_prenodetwo_12_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9176w(0) <= y_prenodetwo_12_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9178w(0) <= y_prenodetwo_12_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9180w(0) <= y_prenodetwo_12_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9182w(0) <= y_prenodetwo_12_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9184w(0) <= y_prenodetwo_12_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9186w(0) <= y_prenodetwo_12_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9335w(0) <= y_prenodetwo_12_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9188w(0) <= y_prenodetwo_12_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9190w(0) <= y_prenodetwo_12_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9192w(0) <= y_prenodetwo_12_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9194w(0) <= y_prenodetwo_12_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9338w(0) <= y_prenodetwo_12_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9341w(0) <= y_prenodetwo_12_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9344w(0) <= y_prenodetwo_12_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9347w(0) <= y_prenodetwo_12_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9350w(0) <= y_prenodetwo_12_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9353w(0) <= y_prenodetwo_12_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9356w(0) <= y_prenodetwo_12_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10130w(0) <= y_prenodetwo_13_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10159w(0) <= y_prenodetwo_13_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10162w(0) <= y_prenodetwo_13_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10165w(0) <= y_prenodetwo_13_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10168w(0) <= y_prenodetwo_13_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10171w(0) <= y_prenodetwo_13_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10174w(0) <= y_prenodetwo_13_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10177w(0) <= y_prenodetwo_13_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10180w(0) <= y_prenodetwo_13_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10183w(0) <= y_prenodetwo_13_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10186w(0) <= y_prenodetwo_13_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10132w(0) <= y_prenodetwo_13_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9973w(0) <= y_prenodetwo_13_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9976w(0) <= y_prenodetwo_13_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9978w(0) <= y_prenodetwo_13_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9980w(0) <= y_prenodetwo_13_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9982w(0) <= y_prenodetwo_13_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9984w(0) <= y_prenodetwo_13_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9986w(0) <= y_prenodetwo_13_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9988w(0) <= y_prenodetwo_13_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9990w(0) <= y_prenodetwo_13_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9992w(0) <= y_prenodetwo_13_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10135w(0) <= y_prenodetwo_13_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9994w(0) <= y_prenodetwo_13_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9996w(0) <= y_prenodetwo_13_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9998w(0) <= y_prenodetwo_13_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10000w(0) <= y_prenodetwo_13_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10138w(0) <= y_prenodetwo_13_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10141w(0) <= y_prenodetwo_13_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10144w(0) <= y_prenodetwo_13_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10147w(0) <= y_prenodetwo_13_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10150w(0) <= y_prenodetwo_13_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10153w(0) <= y_prenodetwo_13_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10156w(0) <= y_prenodetwo_13_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1055w(0) <= y_prenodetwo_2_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1084w(0) <= y_prenodetwo_2_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1087w(0) <= y_prenodetwo_2_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1090w(0) <= y_prenodetwo_2_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1093w(0) <= y_prenodetwo_2_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1096w(0) <= y_prenodetwo_2_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1099w(0) <= y_prenodetwo_2_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1102w(0) <= y_prenodetwo_2_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1105w(0) <= y_prenodetwo_2_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1108w(0) <= y_prenodetwo_2_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1111w(0) <= y_prenodetwo_2_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1057w(0) <= y_prenodetwo_2_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1114w(0) <= y_prenodetwo_2_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1117w(0) <= y_prenodetwo_2_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1120w(0) <= y_prenodetwo_2_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1123w(0) <= y_prenodetwo_2_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1126w(0) <= y_prenodetwo_2_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1129w(0) <= y_prenodetwo_2_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1132w(0) <= y_prenodetwo_2_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1135w(0) <= y_prenodetwo_2_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1138w(0) <= y_prenodetwo_2_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1141w(0) <= y_prenodetwo_2_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1060w(0) <= y_prenodetwo_2_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1144w(0) <= y_prenodetwo_2_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range854w(0) <= y_prenodetwo_2_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range857w(0) <= y_prenodetwo_2_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range859w(0) <= y_prenodetwo_2_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1063w(0) <= y_prenodetwo_2_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1066w(0) <= y_prenodetwo_2_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1069w(0) <= y_prenodetwo_2_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1072w(0) <= y_prenodetwo_2_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1075w(0) <= y_prenodetwo_2_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1078w(0) <= y_prenodetwo_2_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1081w(0) <= y_prenodetwo_2_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1905w(0) <= y_prenodetwo_3_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1934w(0) <= y_prenodetwo_3_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1937w(0) <= y_prenodetwo_3_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1940w(0) <= y_prenodetwo_3_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1943w(0) <= y_prenodetwo_3_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1946w(0) <= y_prenodetwo_3_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1949w(0) <= y_prenodetwo_3_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1952w(0) <= y_prenodetwo_3_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1955w(0) <= y_prenodetwo_3_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1958w(0) <= y_prenodetwo_3_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1961w(0) <= y_prenodetwo_3_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1907w(0) <= y_prenodetwo_3_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1964w(0) <= y_prenodetwo_3_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1967w(0) <= y_prenodetwo_3_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1970w(0) <= y_prenodetwo_3_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1973w(0) <= y_prenodetwo_3_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1976w(0) <= y_prenodetwo_3_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1979w(0) <= y_prenodetwo_3_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1982w(0) <= y_prenodetwo_3_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1985w(0) <= y_prenodetwo_3_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1988w(0) <= y_prenodetwo_3_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1991w(0) <= y_prenodetwo_3_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1910w(0) <= y_prenodetwo_3_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1708w(0) <= y_prenodetwo_3_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1711w(0) <= y_prenodetwo_3_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1713w(0) <= y_prenodetwo_3_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1715w(0) <= y_prenodetwo_3_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1913w(0) <= y_prenodetwo_3_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1916w(0) <= y_prenodetwo_3_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1919w(0) <= y_prenodetwo_3_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1922w(0) <= y_prenodetwo_3_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1925w(0) <= y_prenodetwo_3_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1928w(0) <= y_prenodetwo_3_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1931w(0) <= y_prenodetwo_3_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2750w(0) <= y_prenodetwo_4_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2779w(0) <= y_prenodetwo_4_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2782w(0) <= y_prenodetwo_4_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2785w(0) <= y_prenodetwo_4_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2788w(0) <= y_prenodetwo_4_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2791w(0) <= y_prenodetwo_4_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2794w(0) <= y_prenodetwo_4_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2797w(0) <= y_prenodetwo_4_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2800w(0) <= y_prenodetwo_4_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2803w(0) <= y_prenodetwo_4_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2806w(0) <= y_prenodetwo_4_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2752w(0) <= y_prenodetwo_4_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2809w(0) <= y_prenodetwo_4_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2812w(0) <= y_prenodetwo_4_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2815w(0) <= y_prenodetwo_4_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2818w(0) <= y_prenodetwo_4_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2821w(0) <= y_prenodetwo_4_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2824w(0) <= y_prenodetwo_4_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2827w(0) <= y_prenodetwo_4_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2830w(0) <= y_prenodetwo_4_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2833w(0) <= y_prenodetwo_4_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2557w(0) <= y_prenodetwo_4_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2755w(0) <= y_prenodetwo_4_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2560w(0) <= y_prenodetwo_4_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2562w(0) <= y_prenodetwo_4_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2564w(0) <= y_prenodetwo_4_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2566w(0) <= y_prenodetwo_4_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2758w(0) <= y_prenodetwo_4_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2761w(0) <= y_prenodetwo_4_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2764w(0) <= y_prenodetwo_4_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2767w(0) <= y_prenodetwo_4_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2770w(0) <= y_prenodetwo_4_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2773w(0) <= y_prenodetwo_4_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2776w(0) <= y_prenodetwo_4_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3590w(0) <= y_prenodetwo_5_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3619w(0) <= y_prenodetwo_5_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3622w(0) <= y_prenodetwo_5_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3625w(0) <= y_prenodetwo_5_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3628w(0) <= y_prenodetwo_5_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3631w(0) <= y_prenodetwo_5_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3634w(0) <= y_prenodetwo_5_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3637w(0) <= y_prenodetwo_5_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3640w(0) <= y_prenodetwo_5_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3643w(0) <= y_prenodetwo_5_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3646w(0) <= y_prenodetwo_5_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3592w(0) <= y_prenodetwo_5_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3649w(0) <= y_prenodetwo_5_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3652w(0) <= y_prenodetwo_5_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3655w(0) <= y_prenodetwo_5_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3658w(0) <= y_prenodetwo_5_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3661w(0) <= y_prenodetwo_5_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3664w(0) <= y_prenodetwo_5_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3667w(0) <= y_prenodetwo_5_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3670w(0) <= y_prenodetwo_5_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3401w(0) <= y_prenodetwo_5_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3404w(0) <= y_prenodetwo_5_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3595w(0) <= y_prenodetwo_5_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3406w(0) <= y_prenodetwo_5_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3408w(0) <= y_prenodetwo_5_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3410w(0) <= y_prenodetwo_5_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3412w(0) <= y_prenodetwo_5_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3598w(0) <= y_prenodetwo_5_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3601w(0) <= y_prenodetwo_5_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3604w(0) <= y_prenodetwo_5_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3607w(0) <= y_prenodetwo_5_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3610w(0) <= y_prenodetwo_5_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3613w(0) <= y_prenodetwo_5_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3616w(0) <= y_prenodetwo_5_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4425w(0) <= y_prenodetwo_6_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4454w(0) <= y_prenodetwo_6_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4457w(0) <= y_prenodetwo_6_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4460w(0) <= y_prenodetwo_6_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4463w(0) <= y_prenodetwo_6_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4466w(0) <= y_prenodetwo_6_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4469w(0) <= y_prenodetwo_6_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4472w(0) <= y_prenodetwo_6_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4475w(0) <= y_prenodetwo_6_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4478w(0) <= y_prenodetwo_6_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4481w(0) <= y_prenodetwo_6_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4427w(0) <= y_prenodetwo_6_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4484w(0) <= y_prenodetwo_6_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4487w(0) <= y_prenodetwo_6_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4490w(0) <= y_prenodetwo_6_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4493w(0) <= y_prenodetwo_6_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4496w(0) <= y_prenodetwo_6_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4499w(0) <= y_prenodetwo_6_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4502w(0) <= y_prenodetwo_6_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4240w(0) <= y_prenodetwo_6_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4243w(0) <= y_prenodetwo_6_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4245w(0) <= y_prenodetwo_6_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4430w(0) <= y_prenodetwo_6_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4247w(0) <= y_prenodetwo_6_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4249w(0) <= y_prenodetwo_6_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4251w(0) <= y_prenodetwo_6_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4253w(0) <= y_prenodetwo_6_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4433w(0) <= y_prenodetwo_6_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4436w(0) <= y_prenodetwo_6_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4439w(0) <= y_prenodetwo_6_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4442w(0) <= y_prenodetwo_6_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4445w(0) <= y_prenodetwo_6_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4448w(0) <= y_prenodetwo_6_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4451w(0) <= y_prenodetwo_6_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5255w(0) <= y_prenodetwo_7_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5284w(0) <= y_prenodetwo_7_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5287w(0) <= y_prenodetwo_7_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5290w(0) <= y_prenodetwo_7_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5293w(0) <= y_prenodetwo_7_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5296w(0) <= y_prenodetwo_7_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5299w(0) <= y_prenodetwo_7_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5302w(0) <= y_prenodetwo_7_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5305w(0) <= y_prenodetwo_7_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5308w(0) <= y_prenodetwo_7_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5311w(0) <= y_prenodetwo_7_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5257w(0) <= y_prenodetwo_7_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5314w(0) <= y_prenodetwo_7_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5317w(0) <= y_prenodetwo_7_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5320w(0) <= y_prenodetwo_7_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5323w(0) <= y_prenodetwo_7_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5326w(0) <= y_prenodetwo_7_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5329w(0) <= y_prenodetwo_7_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5074w(0) <= y_prenodetwo_7_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5077w(0) <= y_prenodetwo_7_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5079w(0) <= y_prenodetwo_7_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5081w(0) <= y_prenodetwo_7_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5260w(0) <= y_prenodetwo_7_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5083w(0) <= y_prenodetwo_7_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5085w(0) <= y_prenodetwo_7_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5087w(0) <= y_prenodetwo_7_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5089w(0) <= y_prenodetwo_7_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5263w(0) <= y_prenodetwo_7_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5266w(0) <= y_prenodetwo_7_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5269w(0) <= y_prenodetwo_7_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5272w(0) <= y_prenodetwo_7_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5275w(0) <= y_prenodetwo_7_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5278w(0) <= y_prenodetwo_7_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5281w(0) <= y_prenodetwo_7_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6080w(0) <= y_prenodetwo_8_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6109w(0) <= y_prenodetwo_8_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6112w(0) <= y_prenodetwo_8_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6115w(0) <= y_prenodetwo_8_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6118w(0) <= y_prenodetwo_8_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6121w(0) <= y_prenodetwo_8_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6124w(0) <= y_prenodetwo_8_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6127w(0) <= y_prenodetwo_8_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6130w(0) <= y_prenodetwo_8_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6133w(0) <= y_prenodetwo_8_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6136w(0) <= y_prenodetwo_8_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6082w(0) <= y_prenodetwo_8_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6139w(0) <= y_prenodetwo_8_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6142w(0) <= y_prenodetwo_8_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6145w(0) <= y_prenodetwo_8_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6148w(0) <= y_prenodetwo_8_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6151w(0) <= y_prenodetwo_8_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5903w(0) <= y_prenodetwo_8_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5906w(0) <= y_prenodetwo_8_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5908w(0) <= y_prenodetwo_8_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5910w(0) <= y_prenodetwo_8_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5912w(0) <= y_prenodetwo_8_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6085w(0) <= y_prenodetwo_8_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5914w(0) <= y_prenodetwo_8_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5916w(0) <= y_prenodetwo_8_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5918w(0) <= y_prenodetwo_8_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5920w(0) <= y_prenodetwo_8_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6088w(0) <= y_prenodetwo_8_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6091w(0) <= y_prenodetwo_8_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6094w(0) <= y_prenodetwo_8_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6097w(0) <= y_prenodetwo_8_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6100w(0) <= y_prenodetwo_8_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6103w(0) <= y_prenodetwo_8_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6106w(0) <= y_prenodetwo_8_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6900w(0) <= y_prenodetwo_9_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6929w(0) <= y_prenodetwo_9_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6932w(0) <= y_prenodetwo_9_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6935w(0) <= y_prenodetwo_9_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6938w(0) <= y_prenodetwo_9_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6941w(0) <= y_prenodetwo_9_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6944w(0) <= y_prenodetwo_9_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6947w(0) <= y_prenodetwo_9_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6950w(0) <= y_prenodetwo_9_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6953w(0) <= y_prenodetwo_9_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6956w(0) <= y_prenodetwo_9_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6902w(0) <= y_prenodetwo_9_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6959w(0) <= y_prenodetwo_9_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6962w(0) <= y_prenodetwo_9_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6965w(0) <= y_prenodetwo_9_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6968w(0) <= y_prenodetwo_9_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6727w(0) <= y_prenodetwo_9_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6730w(0) <= y_prenodetwo_9_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6732w(0) <= y_prenodetwo_9_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6734w(0) <= y_prenodetwo_9_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6736w(0) <= y_prenodetwo_9_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6738w(0) <= y_prenodetwo_9_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6905w(0) <= y_prenodetwo_9_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6740w(0) <= y_prenodetwo_9_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6742w(0) <= y_prenodetwo_9_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6744w(0) <= y_prenodetwo_9_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6746w(0) <= y_prenodetwo_9_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6908w(0) <= y_prenodetwo_9_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6911w(0) <= y_prenodetwo_9_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6914w(0) <= y_prenodetwo_9_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6917w(0) <= y_prenodetwo_9_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6920w(0) <= y_prenodetwo_9_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6923w(0) <= y_prenodetwo_9_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6926w(0) <= y_prenodetwo_9_w(9);
	cata_0_cordic_atan :  mysincos_altfp_sincos_cordic_atan_08b
	  PORT MAP ( 
		arctan => wire_cata_0_cordic_atan_arctan,
		indexbit => indexbitff(0)
	  );
	cata_10_cordic_atan :  mysincos_altfp_sincos_cordic_atan_h9b
	  PORT MAP ( 
		arctan => wire_cata_10_cordic_atan_arctan,
		indexbit => indexbitff(10)
	  );
	cata_11_cordic_atan :  mysincos_altfp_sincos_cordic_atan_i9b
	  PORT MAP ( 
		arctan => wire_cata_11_cordic_atan_arctan,
		indexbit => indexbitff(11)
	  );
	cata_12_cordic_atan :  mysincos_altfp_sincos_cordic_atan_j9b
	  PORT MAP ( 
		arctan => wire_cata_12_cordic_atan_arctan,
		indexbit => indexbitff(12)
	  );
	cata_13_cordic_atan :  mysincos_altfp_sincos_cordic_atan_k9b
	  PORT MAP ( 
		arctan => wire_cata_13_cordic_atan_arctan,
		indexbit => indexbitff(13)
	  );
	cata_1_cordic_atan :  mysincos_altfp_sincos_cordic_atan_18b
	  PORT MAP ( 
		arctan => wire_cata_1_cordic_atan_arctan,
		indexbit => indexbitff(1)
	  );
	cata_2_cordic_atan :  mysincos_altfp_sincos_cordic_atan_28b
	  PORT MAP ( 
		arctan => wire_cata_2_cordic_atan_arctan,
		indexbit => indexbitff(2)
	  );
	cata_3_cordic_atan :  mysincos_altfp_sincos_cordic_atan_38b
	  PORT MAP ( 
		arctan => wire_cata_3_cordic_atan_arctan,
		indexbit => indexbitff(3)
	  );
	cata_4_cordic_atan :  mysincos_altfp_sincos_cordic_atan_48b
	  PORT MAP ( 
		arctan => wire_cata_4_cordic_atan_arctan,
		indexbit => indexbitff(4)
	  );
	cata_5_cordic_atan :  mysincos_altfp_sincos_cordic_atan_58b
	  PORT MAP ( 
		arctan => wire_cata_5_cordic_atan_arctan,
		indexbit => indexbitff(5)
	  );
	cata_6_cordic_atan :  mysincos_altfp_sincos_cordic_atan_68b
	  PORT MAP ( 
		arctan => wire_cata_6_cordic_atan_arctan,
		indexbit => indexbitff(6)
	  );
	cata_7_cordic_atan :  mysincos_altfp_sincos_cordic_atan_78b
	  PORT MAP ( 
		arctan => wire_cata_7_cordic_atan_arctan,
		indexbit => indexbitff(7)
	  );
	cata_8_cordic_atan :  mysincos_altfp_sincos_cordic_atan_88b
	  PORT MAP ( 
		arctan => wire_cata_8_cordic_atan_arctan,
		indexbit => indexbitff(8)
	  );
	cata_9_cordic_atan :  mysincos_altfp_sincos_cordic_atan_98b
	  PORT MAP ( 
		arctan => wire_cata_9_cordic_atan_arctan,
		indexbit => indexbitff(9)
	  );
	cxs :  mysincos_altfp_sincos_cordic_start_339
	  PORT MAP ( 
		index => startindex_w,
		value => wire_cxs_value
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cdaff_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cdaff_0 <= delay_input_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cdaff_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cdaff_1 <= cdaff_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cdaff_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cdaff_2 <= cdaff_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN indexbitff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN indexbitff <= ( indexbitff(15 DOWNTO 0) & indexbit);
			END IF;
		END IF;
	END PROCESS;
	wire_indexbitff_w_lg_w_q_range581w681w(0) <= NOT wire_indexbitff_w_q_range581w(0);
	wire_indexbitff_w_lg_w_q_range610w8591w(0) <= NOT wire_indexbitff_w_q_range610w(0);
	wire_indexbitff_w_lg_w_q_range613w9393w(0) <= NOT wire_indexbitff_w_q_range613w(0);
	wire_indexbitff_w_lg_w_q_range616w10190w(0) <= NOT wire_indexbitff_w_q_range616w(0);
	wire_indexbitff_w_lg_w_q_range10749w10754w(0) <= NOT wire_indexbitff_w_q_range10749w(0);
	wire_indexbitff_w_lg_w_q_range583w1148w(0) <= NOT wire_indexbitff_w_q_range583w(0);
	wire_indexbitff_w_lg_w_q_range586w1995w(0) <= NOT wire_indexbitff_w_q_range586w(0);
	wire_indexbitff_w_lg_w_q_range589w2837w(0) <= NOT wire_indexbitff_w_q_range589w(0);
	wire_indexbitff_w_lg_w_q_range592w3674w(0) <= NOT wire_indexbitff_w_q_range592w(0);
	wire_indexbitff_w_lg_w_q_range595w4506w(0) <= NOT wire_indexbitff_w_q_range595w(0);
	wire_indexbitff_w_lg_w_q_range598w5333w(0) <= NOT wire_indexbitff_w_q_range598w(0);
	wire_indexbitff_w_lg_w_q_range601w6155w(0) <= NOT wire_indexbitff_w_q_range601w(0);
	wire_indexbitff_w_lg_w_q_range604w6972w(0) <= NOT wire_indexbitff_w_q_range604w(0);
	wire_indexbitff_w_lg_w_q_range607w7784w(0) <= NOT wire_indexbitff_w_q_range607w(0);
	wire_indexbitff_w_q_range581w(0) <= indexbitff(0);
	wire_indexbitff_w_q_range610w(0) <= indexbitff(10);
	wire_indexbitff_w_q_range613w(0) <= indexbitff(11);
	wire_indexbitff_w_q_range616w(0) <= indexbitff(12);
	wire_indexbitff_w_q_range10749w(0) <= indexbitff(16);
	wire_indexbitff_w_q_range583w(0) <= indexbitff(1);
	wire_indexbitff_w_q_range586w(0) <= indexbitff(2);
	wire_indexbitff_w_q_range589w(0) <= indexbitff(3);
	wire_indexbitff_w_q_range592w(0) <= indexbitff(4);
	wire_indexbitff_w_q_range595w(0) <= indexbitff(5);
	wire_indexbitff_w_q_range598w(0) <= indexbitff(6);
	wire_indexbitff_w_q_range601w(0) <= indexbitff(7);
	wire_indexbitff_w_q_range604w(0) <= indexbitff(8);
	wire_indexbitff_w_q_range607w(0) <= indexbitff(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sincosbitff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN sincosbitff <= ( sincosbitff(15 DOWNTO 0) & sincosbit);
			END IF;
		END IF;
	END PROCESS;
	wire_sincosbitff_w_lg_w_q_range668w10739w(0) <= NOT wire_sincosbitff_w_q_range668w(0);
	wire_sincosbitff_w_lg_w_q_range10746w10747w(0) <= NOT wire_sincosbitff_w_q_range10746w(0);
	wire_sincosbitff_w_q_range668w(0) <= sincosbitff(13);
	wire_sincosbitff_w_q_range10746w(0) <= sincosbitff(16);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sincosff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN sincosff <= wire_sincos_add_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_0 <= x_start_node_w;
			END IF;
		END IF;
	END PROCESS;
	wire_x_pipeff_0_w_lg_w_q_range678w682w(0) <= wire_x_pipeff_0_w_q_range678w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range721w734w(0) <= wire_x_pipeff_0_w_q_range721w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range721w723w(0) <= wire_x_pipeff_0_w_q_range721w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range726w739w(0) <= wire_x_pipeff_0_w_q_range726w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range726w728w(0) <= wire_x_pipeff_0_w_q_range726w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range731w744w(0) <= wire_x_pipeff_0_w_q_range731w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range731w733w(0) <= wire_x_pipeff_0_w_q_range731w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range736w749w(0) <= wire_x_pipeff_0_w_q_range736w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range736w738w(0) <= wire_x_pipeff_0_w_q_range736w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range741w754w(0) <= wire_x_pipeff_0_w_q_range741w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range741w743w(0) <= wire_x_pipeff_0_w_q_range741w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range746w759w(0) <= wire_x_pipeff_0_w_q_range746w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range746w748w(0) <= wire_x_pipeff_0_w_q_range746w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range751w764w(0) <= wire_x_pipeff_0_w_q_range751w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range751w753w(0) <= wire_x_pipeff_0_w_q_range751w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range756w769w(0) <= wire_x_pipeff_0_w_q_range756w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range756w758w(0) <= wire_x_pipeff_0_w_q_range756w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range761w774w(0) <= wire_x_pipeff_0_w_q_range761w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range761w763w(0) <= wire_x_pipeff_0_w_q_range761w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range766w779w(0) <= wire_x_pipeff_0_w_q_range766w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range766w768w(0) <= wire_x_pipeff_0_w_q_range766w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range686w689w(0) <= wire_x_pipeff_0_w_q_range686w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range771w784w(0) <= wire_x_pipeff_0_w_q_range771w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range771w773w(0) <= wire_x_pipeff_0_w_q_range771w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range776w789w(0) <= wire_x_pipeff_0_w_q_range776w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range776w778w(0) <= wire_x_pipeff_0_w_q_range776w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range781w794w(0) <= wire_x_pipeff_0_w_q_range781w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range781w783w(0) <= wire_x_pipeff_0_w_q_range781w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range786w799w(0) <= wire_x_pipeff_0_w_q_range786w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range786w788w(0) <= wire_x_pipeff_0_w_q_range786w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range791w804w(0) <= wire_x_pipeff_0_w_q_range791w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range791w793w(0) <= wire_x_pipeff_0_w_q_range791w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range796w809w(0) <= wire_x_pipeff_0_w_q_range796w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range796w798w(0) <= wire_x_pipeff_0_w_q_range796w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range801w814w(0) <= wire_x_pipeff_0_w_q_range801w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range801w803w(0) <= wire_x_pipeff_0_w_q_range801w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range806w819w(0) <= wire_x_pipeff_0_w_q_range806w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range806w808w(0) <= wire_x_pipeff_0_w_q_range806w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range811w824w(0) <= wire_x_pipeff_0_w_q_range811w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range811w813w(0) <= wire_x_pipeff_0_w_q_range811w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range816w829w(0) <= wire_x_pipeff_0_w_q_range816w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range816w818w(0) <= wire_x_pipeff_0_w_q_range816w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range677w694w(0) <= wire_x_pipeff_0_w_q_range677w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range677w680w(0) <= wire_x_pipeff_0_w_q_range677w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range821w834w(0) <= wire_x_pipeff_0_w_q_range821w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range821w823w(0) <= wire_x_pipeff_0_w_q_range821w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range826w839w(0) <= wire_x_pipeff_0_w_q_range826w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range826w828w(0) <= wire_x_pipeff_0_w_q_range826w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range831w842w(0) <= wire_x_pipeff_0_w_q_range831w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range831w833w(0) <= wire_x_pipeff_0_w_q_range831w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range836w838w(0) <= wire_x_pipeff_0_w_q_range836w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range685w699w(0) <= wire_x_pipeff_0_w_q_range685w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range685w688w(0) <= wire_x_pipeff_0_w_q_range685w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range691w704w(0) <= wire_x_pipeff_0_w_q_range691w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range691w693w(0) <= wire_x_pipeff_0_w_q_range691w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range696w709w(0) <= wire_x_pipeff_0_w_q_range696w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range696w698w(0) <= wire_x_pipeff_0_w_q_range696w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range701w714w(0) <= wire_x_pipeff_0_w_q_range701w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range701w703w(0) <= wire_x_pipeff_0_w_q_range701w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range706w719w(0) <= wire_x_pipeff_0_w_q_range706w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range706w708w(0) <= wire_x_pipeff_0_w_q_range706w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range711w724w(0) <= wire_x_pipeff_0_w_q_range711w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range711w713w(0) <= wire_x_pipeff_0_w_q_range711w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range716w729w(0) <= wire_x_pipeff_0_w_q_range716w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_q_range716w718w(0) <= wire_x_pipeff_0_w_q_range716w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range836w844w(0) <= wire_x_pipeff_0_w_q_range836w(0) AND wire_indexbitff_w_lg_w_q_range581w681w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range678w682w683w(0) <= wire_x_pipeff_0_w_lg_w_q_range678w682w(0) OR wire_x_pipeff_0_w_lg_w_q_range677w680w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range721w734w735w(0) <= wire_x_pipeff_0_w_lg_w_q_range721w734w(0) OR wire_x_pipeff_0_w_lg_w_q_range731w733w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range726w739w740w(0) <= wire_x_pipeff_0_w_lg_w_q_range726w739w(0) OR wire_x_pipeff_0_w_lg_w_q_range736w738w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range731w744w745w(0) <= wire_x_pipeff_0_w_lg_w_q_range731w744w(0) OR wire_x_pipeff_0_w_lg_w_q_range741w743w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range736w749w750w(0) <= wire_x_pipeff_0_w_lg_w_q_range736w749w(0) OR wire_x_pipeff_0_w_lg_w_q_range746w748w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range741w754w755w(0) <= wire_x_pipeff_0_w_lg_w_q_range741w754w(0) OR wire_x_pipeff_0_w_lg_w_q_range751w753w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range746w759w760w(0) <= wire_x_pipeff_0_w_lg_w_q_range746w759w(0) OR wire_x_pipeff_0_w_lg_w_q_range756w758w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range751w764w765w(0) <= wire_x_pipeff_0_w_lg_w_q_range751w764w(0) OR wire_x_pipeff_0_w_lg_w_q_range761w763w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range756w769w770w(0) <= wire_x_pipeff_0_w_lg_w_q_range756w769w(0) OR wire_x_pipeff_0_w_lg_w_q_range766w768w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range761w774w775w(0) <= wire_x_pipeff_0_w_lg_w_q_range761w774w(0) OR wire_x_pipeff_0_w_lg_w_q_range771w773w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range766w779w780w(0) <= wire_x_pipeff_0_w_lg_w_q_range766w779w(0) OR wire_x_pipeff_0_w_lg_w_q_range776w778w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range686w689w690w(0) <= wire_x_pipeff_0_w_lg_w_q_range686w689w(0) OR wire_x_pipeff_0_w_lg_w_q_range685w688w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range771w784w785w(0) <= wire_x_pipeff_0_w_lg_w_q_range771w784w(0) OR wire_x_pipeff_0_w_lg_w_q_range781w783w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range776w789w790w(0) <= wire_x_pipeff_0_w_lg_w_q_range776w789w(0) OR wire_x_pipeff_0_w_lg_w_q_range786w788w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range781w794w795w(0) <= wire_x_pipeff_0_w_lg_w_q_range781w794w(0) OR wire_x_pipeff_0_w_lg_w_q_range791w793w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range786w799w800w(0) <= wire_x_pipeff_0_w_lg_w_q_range786w799w(0) OR wire_x_pipeff_0_w_lg_w_q_range796w798w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range791w804w805w(0) <= wire_x_pipeff_0_w_lg_w_q_range791w804w(0) OR wire_x_pipeff_0_w_lg_w_q_range801w803w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range796w809w810w(0) <= wire_x_pipeff_0_w_lg_w_q_range796w809w(0) OR wire_x_pipeff_0_w_lg_w_q_range806w808w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range801w814w815w(0) <= wire_x_pipeff_0_w_lg_w_q_range801w814w(0) OR wire_x_pipeff_0_w_lg_w_q_range811w813w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range806w819w820w(0) <= wire_x_pipeff_0_w_lg_w_q_range806w819w(0) OR wire_x_pipeff_0_w_lg_w_q_range816w818w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range811w824w825w(0) <= wire_x_pipeff_0_w_lg_w_q_range811w824w(0) OR wire_x_pipeff_0_w_lg_w_q_range821w823w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range816w829w830w(0) <= wire_x_pipeff_0_w_lg_w_q_range816w829w(0) OR wire_x_pipeff_0_w_lg_w_q_range826w828w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range677w694w695w(0) <= wire_x_pipeff_0_w_lg_w_q_range677w694w(0) OR wire_x_pipeff_0_w_lg_w_q_range691w693w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range821w834w835w(0) <= wire_x_pipeff_0_w_lg_w_q_range821w834w(0) OR wire_x_pipeff_0_w_lg_w_q_range831w833w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range826w839w840w(0) <= wire_x_pipeff_0_w_lg_w_q_range826w839w(0) OR wire_x_pipeff_0_w_lg_w_q_range836w838w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range685w699w700w(0) <= wire_x_pipeff_0_w_lg_w_q_range685w699w(0) OR wire_x_pipeff_0_w_lg_w_q_range696w698w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range691w704w705w(0) <= wire_x_pipeff_0_w_lg_w_q_range691w704w(0) OR wire_x_pipeff_0_w_lg_w_q_range701w703w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range696w709w710w(0) <= wire_x_pipeff_0_w_lg_w_q_range696w709w(0) OR wire_x_pipeff_0_w_lg_w_q_range706w708w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range701w714w715w(0) <= wire_x_pipeff_0_w_lg_w_q_range701w714w(0) OR wire_x_pipeff_0_w_lg_w_q_range711w713w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range706w719w720w(0) <= wire_x_pipeff_0_w_lg_w_q_range706w719w(0) OR wire_x_pipeff_0_w_lg_w_q_range716w718w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range711w724w725w(0) <= wire_x_pipeff_0_w_lg_w_q_range711w724w(0) OR wire_x_pipeff_0_w_lg_w_q_range721w723w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range716w729w730w(0) <= wire_x_pipeff_0_w_lg_w_q_range716w729w(0) OR wire_x_pipeff_0_w_lg_w_q_range726w728w(0);
	wire_x_pipeff_0_w_q_range678w(0) <= x_pipeff_0(0);
	wire_x_pipeff_0_w_q_range721w(0) <= x_pipeff_0(10);
	wire_x_pipeff_0_w_q_range726w(0) <= x_pipeff_0(11);
	wire_x_pipeff_0_w_q_range731w(0) <= x_pipeff_0(12);
	wire_x_pipeff_0_w_q_range736w(0) <= x_pipeff_0(13);
	wire_x_pipeff_0_w_q_range741w(0) <= x_pipeff_0(14);
	wire_x_pipeff_0_w_q_range746w(0) <= x_pipeff_0(15);
	wire_x_pipeff_0_w_q_range751w(0) <= x_pipeff_0(16);
	wire_x_pipeff_0_w_q_range756w(0) <= x_pipeff_0(17);
	wire_x_pipeff_0_w_q_range761w(0) <= x_pipeff_0(18);
	wire_x_pipeff_0_w_q_range766w(0) <= x_pipeff_0(19);
	wire_x_pipeff_0_w_q_range686w(0) <= x_pipeff_0(1);
	wire_x_pipeff_0_w_q_range771w(0) <= x_pipeff_0(20);
	wire_x_pipeff_0_w_q_range776w(0) <= x_pipeff_0(21);
	wire_x_pipeff_0_w_q_range781w(0) <= x_pipeff_0(22);
	wire_x_pipeff_0_w_q_range786w(0) <= x_pipeff_0(23);
	wire_x_pipeff_0_w_q_range791w(0) <= x_pipeff_0(24);
	wire_x_pipeff_0_w_q_range796w(0) <= x_pipeff_0(25);
	wire_x_pipeff_0_w_q_range801w(0) <= x_pipeff_0(26);
	wire_x_pipeff_0_w_q_range806w(0) <= x_pipeff_0(27);
	wire_x_pipeff_0_w_q_range811w(0) <= x_pipeff_0(28);
	wire_x_pipeff_0_w_q_range816w(0) <= x_pipeff_0(29);
	wire_x_pipeff_0_w_q_range677w(0) <= x_pipeff_0(2);
	wire_x_pipeff_0_w_q_range821w(0) <= x_pipeff_0(30);
	wire_x_pipeff_0_w_q_range826w(0) <= x_pipeff_0(31);
	wire_x_pipeff_0_w_q_range831w(0) <= x_pipeff_0(32);
	wire_x_pipeff_0_w_q_range836w(0) <= x_pipeff_0(33);
	wire_x_pipeff_0_w_q_range685w(0) <= x_pipeff_0(3);
	wire_x_pipeff_0_w_q_range691w(0) <= x_pipeff_0(4);
	wire_x_pipeff_0_w_q_range696w(0) <= x_pipeff_0(5);
	wire_x_pipeff_0_w_q_range701w(0) <= x_pipeff_0(6);
	wire_x_pipeff_0_w_q_range706w(0) <= x_pipeff_0(7);
	wire_x_pipeff_0_w_q_range711w(0) <= x_pipeff_0(8);
	wire_x_pipeff_0_w_q_range716w(0) <= x_pipeff_0(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_1 <= x_pipeff_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_10 <= x_pipenode_10_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_11 <= x_pipenode_11_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_12 <= x_pipenode_12_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_13 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_13 <= x_pipenode_13_w;
			END IF;
		END IF;
	END PROCESS;
	loop32 : FOR i IN 0 TO 33 GENERATE 
		wire_x_pipeff_13_w_lg_q10744w(i) <= x_pipeff_13(i) AND wire_sincosbitff_w_lg_w_q_range668w10739w(0);
	END GENERATE loop32;
	loop33 : FOR i IN 0 TO 33 GENERATE 
		wire_x_pipeff_13_w_lg_q10741w(i) <= x_pipeff_13(i) AND wire_sincosbitff_w_q_range668w(0);
	END GENERATE loop33;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_2 <= x_pipenode_2_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_3 <= x_pipenode_3_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_4 <= x_pipenode_4_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_5 <= x_pipenode_5_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_6 <= x_pipenode_6_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_7 <= x_pipenode_7_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_8 <= x_pipenode_8_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_9 <= x_pipenode_9_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(0) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(0) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(1) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(1) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(2) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(2) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(3) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(3) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(4) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(4) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(5) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(5) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(6) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(6) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(7) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(7) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(8) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(8) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(9) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(9) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(10) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(10) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(11) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(11) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(12) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(12) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(13) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(13) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(14) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(14) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(15) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(15) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(16) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(16) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(17) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(17) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(18) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(18) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(19) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(19) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(20) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(20) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(21) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(21) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(22) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(22) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(23) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(23) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(24) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(24) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(25) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(25) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(26) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(26) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(27) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(27) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(28) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(28) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(29) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(29) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(30) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(30) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(31) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(31) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(32) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(32) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(33) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(33) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_1 <= wire_y_pipeff1_add_result;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_1_w_lg_w_q_range913w915w(0) <= NOT wire_y_pipeff_1_w_q_range913w(0);
	wire_y_pipeff_1_w_lg_w_q_range919w921w(0) <= NOT wire_y_pipeff_1_w_q_range919w(0);
	wire_y_pipeff_1_w_lg_w_q_range925w927w(0) <= NOT wire_y_pipeff_1_w_q_range925w(0);
	wire_y_pipeff_1_w_lg_w_q_range931w933w(0) <= NOT wire_y_pipeff_1_w_q_range931w(0);
	wire_y_pipeff_1_w_lg_w_q_range937w939w(0) <= NOT wire_y_pipeff_1_w_q_range937w(0);
	wire_y_pipeff_1_w_lg_w_q_range943w945w(0) <= NOT wire_y_pipeff_1_w_q_range943w(0);
	wire_y_pipeff_1_w_lg_w_q_range949w951w(0) <= NOT wire_y_pipeff_1_w_q_range949w(0);
	wire_y_pipeff_1_w_lg_w_q_range955w957w(0) <= NOT wire_y_pipeff_1_w_q_range955w(0);
	wire_y_pipeff_1_w_lg_w_q_range961w963w(0) <= NOT wire_y_pipeff_1_w_q_range961w(0);
	wire_y_pipeff_1_w_lg_w_q_range967w969w(0) <= NOT wire_y_pipeff_1_w_q_range967w(0);
	wire_y_pipeff_1_w_lg_w_q_range860w862w(0) <= NOT wire_y_pipeff_1_w_q_range860w(0);
	wire_y_pipeff_1_w_lg_w_q_range973w975w(0) <= NOT wire_y_pipeff_1_w_q_range973w(0);
	wire_y_pipeff_1_w_lg_w_q_range979w981w(0) <= NOT wire_y_pipeff_1_w_q_range979w(0);
	wire_y_pipeff_1_w_lg_w_q_range985w987w(0) <= NOT wire_y_pipeff_1_w_q_range985w(0);
	wire_y_pipeff_1_w_lg_w_q_range991w993w(0) <= NOT wire_y_pipeff_1_w_q_range991w(0);
	wire_y_pipeff_1_w_lg_w_q_range997w999w(0) <= NOT wire_y_pipeff_1_w_q_range997w(0);
	wire_y_pipeff_1_w_lg_w_q_range1003w1005w(0) <= NOT wire_y_pipeff_1_w_q_range1003w(0);
	wire_y_pipeff_1_w_lg_w_q_range1009w1011w(0) <= NOT wire_y_pipeff_1_w_q_range1009w(0);
	wire_y_pipeff_1_w_lg_w_q_range1015w1017w(0) <= NOT wire_y_pipeff_1_w_q_range1015w(0);
	wire_y_pipeff_1_w_lg_w_q_range1021w1023w(0) <= NOT wire_y_pipeff_1_w_q_range1021w(0);
	wire_y_pipeff_1_w_lg_w_q_range1027w1029w(0) <= NOT wire_y_pipeff_1_w_q_range1027w(0);
	wire_y_pipeff_1_w_lg_w_q_range865w867w(0) <= NOT wire_y_pipeff_1_w_q_range865w(0);
	wire_y_pipeff_1_w_lg_w_q_range1033w1035w(0) <= NOT wire_y_pipeff_1_w_q_range1033w(0);
	wire_y_pipeff_1_w_lg_w_q_range1039w1041w(0) <= NOT wire_y_pipeff_1_w_q_range1039w(0);
	wire_y_pipeff_1_w_lg_w_q_range1045w1047w(0) <= NOT wire_y_pipeff_1_w_q_range1045w(0);
	wire_y_pipeff_1_w_lg_w_q_range845w847w(0) <= NOT wire_y_pipeff_1_w_q_range845w(0);
	wire_y_pipeff_1_w_lg_w_q_range871w873w(0) <= NOT wire_y_pipeff_1_w_q_range871w(0);
	wire_y_pipeff_1_w_lg_w_q_range877w879w(0) <= NOT wire_y_pipeff_1_w_q_range877w(0);
	wire_y_pipeff_1_w_lg_w_q_range883w885w(0) <= NOT wire_y_pipeff_1_w_q_range883w(0);
	wire_y_pipeff_1_w_lg_w_q_range889w891w(0) <= NOT wire_y_pipeff_1_w_q_range889w(0);
	wire_y_pipeff_1_w_lg_w_q_range895w897w(0) <= NOT wire_y_pipeff_1_w_q_range895w(0);
	wire_y_pipeff_1_w_lg_w_q_range901w903w(0) <= NOT wire_y_pipeff_1_w_q_range901w(0);
	wire_y_pipeff_1_w_lg_w_q_range907w909w(0) <= NOT wire_y_pipeff_1_w_q_range907w(0);
	wire_y_pipeff_1_w_q_range913w(0) <= y_pipeff_1(10);
	wire_y_pipeff_1_w_q_range919w(0) <= y_pipeff_1(11);
	wire_y_pipeff_1_w_q_range925w(0) <= y_pipeff_1(12);
	wire_y_pipeff_1_w_q_range931w(0) <= y_pipeff_1(13);
	wire_y_pipeff_1_w_q_range937w(0) <= y_pipeff_1(14);
	wire_y_pipeff_1_w_q_range943w(0) <= y_pipeff_1(15);
	wire_y_pipeff_1_w_q_range949w(0) <= y_pipeff_1(16);
	wire_y_pipeff_1_w_q_range955w(0) <= y_pipeff_1(17);
	wire_y_pipeff_1_w_q_range961w(0) <= y_pipeff_1(18);
	wire_y_pipeff_1_w_q_range967w(0) <= y_pipeff_1(19);
	wire_y_pipeff_1_w_q_range860w(0) <= y_pipeff_1(1);
	wire_y_pipeff_1_w_q_range973w(0) <= y_pipeff_1(20);
	wire_y_pipeff_1_w_q_range979w(0) <= y_pipeff_1(21);
	wire_y_pipeff_1_w_q_range985w(0) <= y_pipeff_1(22);
	wire_y_pipeff_1_w_q_range991w(0) <= y_pipeff_1(23);
	wire_y_pipeff_1_w_q_range997w(0) <= y_pipeff_1(24);
	wire_y_pipeff_1_w_q_range1003w(0) <= y_pipeff_1(25);
	wire_y_pipeff_1_w_q_range1009w(0) <= y_pipeff_1(26);
	wire_y_pipeff_1_w_q_range1015w(0) <= y_pipeff_1(27);
	wire_y_pipeff_1_w_q_range1021w(0) <= y_pipeff_1(28);
	wire_y_pipeff_1_w_q_range1027w(0) <= y_pipeff_1(29);
	wire_y_pipeff_1_w_q_range865w(0) <= y_pipeff_1(2);
	wire_y_pipeff_1_w_q_range1033w(0) <= y_pipeff_1(30);
	wire_y_pipeff_1_w_q_range1039w(0) <= y_pipeff_1(31);
	wire_y_pipeff_1_w_q_range1045w(0) <= y_pipeff_1(32);
	wire_y_pipeff_1_w_q_range845w(0) <= y_pipeff_1(33);
	wire_y_pipeff_1_w_q_range871w(0) <= y_pipeff_1(3);
	wire_y_pipeff_1_w_q_range877w(0) <= y_pipeff_1(4);
	wire_y_pipeff_1_w_q_range883w(0) <= y_pipeff_1(5);
	wire_y_pipeff_1_w_q_range889w(0) <= y_pipeff_1(6);
	wire_y_pipeff_1_w_q_range895w(0) <= y_pipeff_1(7);
	wire_y_pipeff_1_w_q_range901w(0) <= y_pipeff_1(8);
	wire_y_pipeff_1_w_q_range907w(0) <= y_pipeff_1(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_10 <= y_pipenode_10_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_10_w_lg_w_q_range8384w8386w(0) <= NOT wire_y_pipeff_10_w_q_range8384w(0);
	wire_y_pipeff_10_w_lg_w_q_range8389w8391w(0) <= NOT wire_y_pipeff_10_w_q_range8389w(0);
	wire_y_pipeff_10_w_lg_w_q_range8395w8397w(0) <= NOT wire_y_pipeff_10_w_q_range8395w(0);
	wire_y_pipeff_10_w_lg_w_q_range8401w8403w(0) <= NOT wire_y_pipeff_10_w_q_range8401w(0);
	wire_y_pipeff_10_w_lg_w_q_range8407w8409w(0) <= NOT wire_y_pipeff_10_w_q_range8407w(0);
	wire_y_pipeff_10_w_lg_w_q_range8413w8415w(0) <= NOT wire_y_pipeff_10_w_q_range8413w(0);
	wire_y_pipeff_10_w_lg_w_q_range8419w8421w(0) <= NOT wire_y_pipeff_10_w_q_range8419w(0);
	wire_y_pipeff_10_w_lg_w_q_range8425w8427w(0) <= NOT wire_y_pipeff_10_w_q_range8425w(0);
	wire_y_pipeff_10_w_lg_w_q_range8431w8433w(0) <= NOT wire_y_pipeff_10_w_q_range8431w(0);
	wire_y_pipeff_10_w_lg_w_q_range8437w8439w(0) <= NOT wire_y_pipeff_10_w_q_range8437w(0);
	wire_y_pipeff_10_w_lg_w_q_range8443w8445w(0) <= NOT wire_y_pipeff_10_w_q_range8443w(0);
	wire_y_pipeff_10_w_lg_w_q_range8449w8451w(0) <= NOT wire_y_pipeff_10_w_q_range8449w(0);
	wire_y_pipeff_10_w_lg_w_q_range8455w8457w(0) <= NOT wire_y_pipeff_10_w_q_range8455w(0);
	wire_y_pipeff_10_w_lg_w_q_range8461w8463w(0) <= NOT wire_y_pipeff_10_w_q_range8461w(0);
	wire_y_pipeff_10_w_lg_w_q_range8467w8469w(0) <= NOT wire_y_pipeff_10_w_q_range8467w(0);
	wire_y_pipeff_10_w_lg_w_q_range8473w8475w(0) <= NOT wire_y_pipeff_10_w_q_range8473w(0);
	wire_y_pipeff_10_w_lg_w_q_range8479w8481w(0) <= NOT wire_y_pipeff_10_w_q_range8479w(0);
	wire_y_pipeff_10_w_lg_w_q_range8485w8487w(0) <= NOT wire_y_pipeff_10_w_q_range8485w(0);
	wire_y_pipeff_10_w_lg_w_q_range8491w8493w(0) <= NOT wire_y_pipeff_10_w_q_range8491w(0);
	wire_y_pipeff_10_w_lg_w_q_range8497w8499w(0) <= NOT wire_y_pipeff_10_w_q_range8497w(0);
	wire_y_pipeff_10_w_lg_w_q_range8503w8505w(0) <= NOT wire_y_pipeff_10_w_q_range8503w(0);
	wire_y_pipeff_10_w_lg_w_q_range8509w8511w(0) <= NOT wire_y_pipeff_10_w_q_range8509w(0);
	wire_y_pipeff_10_w_lg_w_q_range8515w8517w(0) <= NOT wire_y_pipeff_10_w_q_range8515w(0);
	wire_y_pipeff_10_w_lg_w_q_range8333w8335w(0) <= NOT wire_y_pipeff_10_w_q_range8333w(0);
	wire_y_pipeff_10_w_q_range8384w(0) <= y_pipeff_10(10);
	wire_y_pipeff_10_w_q_range8389w(0) <= y_pipeff_10(11);
	wire_y_pipeff_10_w_q_range8395w(0) <= y_pipeff_10(12);
	wire_y_pipeff_10_w_q_range8401w(0) <= y_pipeff_10(13);
	wire_y_pipeff_10_w_q_range8407w(0) <= y_pipeff_10(14);
	wire_y_pipeff_10_w_q_range8413w(0) <= y_pipeff_10(15);
	wire_y_pipeff_10_w_q_range8419w(0) <= y_pipeff_10(16);
	wire_y_pipeff_10_w_q_range8425w(0) <= y_pipeff_10(17);
	wire_y_pipeff_10_w_q_range8431w(0) <= y_pipeff_10(18);
	wire_y_pipeff_10_w_q_range8437w(0) <= y_pipeff_10(19);
	wire_y_pipeff_10_w_q_range8443w(0) <= y_pipeff_10(20);
	wire_y_pipeff_10_w_q_range8449w(0) <= y_pipeff_10(21);
	wire_y_pipeff_10_w_q_range8455w(0) <= y_pipeff_10(22);
	wire_y_pipeff_10_w_q_range8461w(0) <= y_pipeff_10(23);
	wire_y_pipeff_10_w_q_range8467w(0) <= y_pipeff_10(24);
	wire_y_pipeff_10_w_q_range8473w(0) <= y_pipeff_10(25);
	wire_y_pipeff_10_w_q_range8479w(0) <= y_pipeff_10(26);
	wire_y_pipeff_10_w_q_range8485w(0) <= y_pipeff_10(27);
	wire_y_pipeff_10_w_q_range8491w(0) <= y_pipeff_10(28);
	wire_y_pipeff_10_w_q_range8497w(0) <= y_pipeff_10(29);
	wire_y_pipeff_10_w_q_range8503w(0) <= y_pipeff_10(30);
	wire_y_pipeff_10_w_q_range8509w(0) <= y_pipeff_10(31);
	wire_y_pipeff_10_w_q_range8515w(0) <= y_pipeff_10(32);
	wire_y_pipeff_10_w_q_range8333w(0) <= y_pipeff_10(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_11 <= y_pipenode_11_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_11_w_lg_w_q_range9195w9197w(0) <= NOT wire_y_pipeff_11_w_q_range9195w(0);
	wire_y_pipeff_11_w_lg_w_q_range9200w9202w(0) <= NOT wire_y_pipeff_11_w_q_range9200w(0);
	wire_y_pipeff_11_w_lg_w_q_range9206w9208w(0) <= NOT wire_y_pipeff_11_w_q_range9206w(0);
	wire_y_pipeff_11_w_lg_w_q_range9212w9214w(0) <= NOT wire_y_pipeff_11_w_q_range9212w(0);
	wire_y_pipeff_11_w_lg_w_q_range9218w9220w(0) <= NOT wire_y_pipeff_11_w_q_range9218w(0);
	wire_y_pipeff_11_w_lg_w_q_range9224w9226w(0) <= NOT wire_y_pipeff_11_w_q_range9224w(0);
	wire_y_pipeff_11_w_lg_w_q_range9230w9232w(0) <= NOT wire_y_pipeff_11_w_q_range9230w(0);
	wire_y_pipeff_11_w_lg_w_q_range9236w9238w(0) <= NOT wire_y_pipeff_11_w_q_range9236w(0);
	wire_y_pipeff_11_w_lg_w_q_range9242w9244w(0) <= NOT wire_y_pipeff_11_w_q_range9242w(0);
	wire_y_pipeff_11_w_lg_w_q_range9248w9250w(0) <= NOT wire_y_pipeff_11_w_q_range9248w(0);
	wire_y_pipeff_11_w_lg_w_q_range9254w9256w(0) <= NOT wire_y_pipeff_11_w_q_range9254w(0);
	wire_y_pipeff_11_w_lg_w_q_range9260w9262w(0) <= NOT wire_y_pipeff_11_w_q_range9260w(0);
	wire_y_pipeff_11_w_lg_w_q_range9266w9268w(0) <= NOT wire_y_pipeff_11_w_q_range9266w(0);
	wire_y_pipeff_11_w_lg_w_q_range9272w9274w(0) <= NOT wire_y_pipeff_11_w_q_range9272w(0);
	wire_y_pipeff_11_w_lg_w_q_range9278w9280w(0) <= NOT wire_y_pipeff_11_w_q_range9278w(0);
	wire_y_pipeff_11_w_lg_w_q_range9284w9286w(0) <= NOT wire_y_pipeff_11_w_q_range9284w(0);
	wire_y_pipeff_11_w_lg_w_q_range9290w9292w(0) <= NOT wire_y_pipeff_11_w_q_range9290w(0);
	wire_y_pipeff_11_w_lg_w_q_range9296w9298w(0) <= NOT wire_y_pipeff_11_w_q_range9296w(0);
	wire_y_pipeff_11_w_lg_w_q_range9302w9304w(0) <= NOT wire_y_pipeff_11_w_q_range9302w(0);
	wire_y_pipeff_11_w_lg_w_q_range9308w9310w(0) <= NOT wire_y_pipeff_11_w_q_range9308w(0);
	wire_y_pipeff_11_w_lg_w_q_range9314w9316w(0) <= NOT wire_y_pipeff_11_w_q_range9314w(0);
	wire_y_pipeff_11_w_lg_w_q_range9320w9322w(0) <= NOT wire_y_pipeff_11_w_q_range9320w(0);
	wire_y_pipeff_11_w_lg_w_q_range9140w9142w(0) <= NOT wire_y_pipeff_11_w_q_range9140w(0);
	wire_y_pipeff_11_w_q_range9195w(0) <= y_pipeff_11(11);
	wire_y_pipeff_11_w_q_range9200w(0) <= y_pipeff_11(12);
	wire_y_pipeff_11_w_q_range9206w(0) <= y_pipeff_11(13);
	wire_y_pipeff_11_w_q_range9212w(0) <= y_pipeff_11(14);
	wire_y_pipeff_11_w_q_range9218w(0) <= y_pipeff_11(15);
	wire_y_pipeff_11_w_q_range9224w(0) <= y_pipeff_11(16);
	wire_y_pipeff_11_w_q_range9230w(0) <= y_pipeff_11(17);
	wire_y_pipeff_11_w_q_range9236w(0) <= y_pipeff_11(18);
	wire_y_pipeff_11_w_q_range9242w(0) <= y_pipeff_11(19);
	wire_y_pipeff_11_w_q_range9248w(0) <= y_pipeff_11(20);
	wire_y_pipeff_11_w_q_range9254w(0) <= y_pipeff_11(21);
	wire_y_pipeff_11_w_q_range9260w(0) <= y_pipeff_11(22);
	wire_y_pipeff_11_w_q_range9266w(0) <= y_pipeff_11(23);
	wire_y_pipeff_11_w_q_range9272w(0) <= y_pipeff_11(24);
	wire_y_pipeff_11_w_q_range9278w(0) <= y_pipeff_11(25);
	wire_y_pipeff_11_w_q_range9284w(0) <= y_pipeff_11(26);
	wire_y_pipeff_11_w_q_range9290w(0) <= y_pipeff_11(27);
	wire_y_pipeff_11_w_q_range9296w(0) <= y_pipeff_11(28);
	wire_y_pipeff_11_w_q_range9302w(0) <= y_pipeff_11(29);
	wire_y_pipeff_11_w_q_range9308w(0) <= y_pipeff_11(30);
	wire_y_pipeff_11_w_q_range9314w(0) <= y_pipeff_11(31);
	wire_y_pipeff_11_w_q_range9320w(0) <= y_pipeff_11(32);
	wire_y_pipeff_11_w_q_range9140w(0) <= y_pipeff_11(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_12 <= y_pipenode_12_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_12_w_lg_w_q_range10001w10003w(0) <= NOT wire_y_pipeff_12_w_q_range10001w(0);
	wire_y_pipeff_12_w_lg_w_q_range10006w10008w(0) <= NOT wire_y_pipeff_12_w_q_range10006w(0);
	wire_y_pipeff_12_w_lg_w_q_range10012w10014w(0) <= NOT wire_y_pipeff_12_w_q_range10012w(0);
	wire_y_pipeff_12_w_lg_w_q_range10018w10020w(0) <= NOT wire_y_pipeff_12_w_q_range10018w(0);
	wire_y_pipeff_12_w_lg_w_q_range10024w10026w(0) <= NOT wire_y_pipeff_12_w_q_range10024w(0);
	wire_y_pipeff_12_w_lg_w_q_range10030w10032w(0) <= NOT wire_y_pipeff_12_w_q_range10030w(0);
	wire_y_pipeff_12_w_lg_w_q_range10036w10038w(0) <= NOT wire_y_pipeff_12_w_q_range10036w(0);
	wire_y_pipeff_12_w_lg_w_q_range10042w10044w(0) <= NOT wire_y_pipeff_12_w_q_range10042w(0);
	wire_y_pipeff_12_w_lg_w_q_range10048w10050w(0) <= NOT wire_y_pipeff_12_w_q_range10048w(0);
	wire_y_pipeff_12_w_lg_w_q_range10054w10056w(0) <= NOT wire_y_pipeff_12_w_q_range10054w(0);
	wire_y_pipeff_12_w_lg_w_q_range10060w10062w(0) <= NOT wire_y_pipeff_12_w_q_range10060w(0);
	wire_y_pipeff_12_w_lg_w_q_range10066w10068w(0) <= NOT wire_y_pipeff_12_w_q_range10066w(0);
	wire_y_pipeff_12_w_lg_w_q_range10072w10074w(0) <= NOT wire_y_pipeff_12_w_q_range10072w(0);
	wire_y_pipeff_12_w_lg_w_q_range10078w10080w(0) <= NOT wire_y_pipeff_12_w_q_range10078w(0);
	wire_y_pipeff_12_w_lg_w_q_range10084w10086w(0) <= NOT wire_y_pipeff_12_w_q_range10084w(0);
	wire_y_pipeff_12_w_lg_w_q_range10090w10092w(0) <= NOT wire_y_pipeff_12_w_q_range10090w(0);
	wire_y_pipeff_12_w_lg_w_q_range10096w10098w(0) <= NOT wire_y_pipeff_12_w_q_range10096w(0);
	wire_y_pipeff_12_w_lg_w_q_range10102w10104w(0) <= NOT wire_y_pipeff_12_w_q_range10102w(0);
	wire_y_pipeff_12_w_lg_w_q_range10108w10110w(0) <= NOT wire_y_pipeff_12_w_q_range10108w(0);
	wire_y_pipeff_12_w_lg_w_q_range10114w10116w(0) <= NOT wire_y_pipeff_12_w_q_range10114w(0);
	wire_y_pipeff_12_w_lg_w_q_range10120w10122w(0) <= NOT wire_y_pipeff_12_w_q_range10120w(0);
	wire_y_pipeff_12_w_lg_w_q_range9942w9944w(0) <= NOT wire_y_pipeff_12_w_q_range9942w(0);
	wire_y_pipeff_12_w_q_range10001w(0) <= y_pipeff_12(12);
	wire_y_pipeff_12_w_q_range10006w(0) <= y_pipeff_12(13);
	wire_y_pipeff_12_w_q_range10012w(0) <= y_pipeff_12(14);
	wire_y_pipeff_12_w_q_range10018w(0) <= y_pipeff_12(15);
	wire_y_pipeff_12_w_q_range10024w(0) <= y_pipeff_12(16);
	wire_y_pipeff_12_w_q_range10030w(0) <= y_pipeff_12(17);
	wire_y_pipeff_12_w_q_range10036w(0) <= y_pipeff_12(18);
	wire_y_pipeff_12_w_q_range10042w(0) <= y_pipeff_12(19);
	wire_y_pipeff_12_w_q_range10048w(0) <= y_pipeff_12(20);
	wire_y_pipeff_12_w_q_range10054w(0) <= y_pipeff_12(21);
	wire_y_pipeff_12_w_q_range10060w(0) <= y_pipeff_12(22);
	wire_y_pipeff_12_w_q_range10066w(0) <= y_pipeff_12(23);
	wire_y_pipeff_12_w_q_range10072w(0) <= y_pipeff_12(24);
	wire_y_pipeff_12_w_q_range10078w(0) <= y_pipeff_12(25);
	wire_y_pipeff_12_w_q_range10084w(0) <= y_pipeff_12(26);
	wire_y_pipeff_12_w_q_range10090w(0) <= y_pipeff_12(27);
	wire_y_pipeff_12_w_q_range10096w(0) <= y_pipeff_12(28);
	wire_y_pipeff_12_w_q_range10102w(0) <= y_pipeff_12(29);
	wire_y_pipeff_12_w_q_range10108w(0) <= y_pipeff_12(30);
	wire_y_pipeff_12_w_q_range10114w(0) <= y_pipeff_12(31);
	wire_y_pipeff_12_w_q_range10120w(0) <= y_pipeff_12(32);
	wire_y_pipeff_12_w_q_range9942w(0) <= y_pipeff_12(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_13 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_13 <= y_pipenode_13_w;
			END IF;
		END IF;
	END PROCESS;
	loop34 : FOR i IN 0 TO 33 GENERATE 
		wire_y_pipeff_13_w_lg_q10740w(i) <= y_pipeff_13(i) AND wire_sincosbitff_w_lg_w_q_range668w10739w(0);
	END GENERATE loop34;
	loop35 : FOR i IN 0 TO 33 GENERATE 
		wire_y_pipeff_13_w_lg_q10743w(i) <= y_pipeff_13(i) AND wire_sincosbitff_w_q_range668w(0);
	END GENERATE loop35;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_2 <= y_pipenode_2_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_2_w_lg_w_q_range1763w1765w(0) <= NOT wire_y_pipeff_2_w_q_range1763w(0);
	wire_y_pipeff_2_w_lg_w_q_range1769w1771w(0) <= NOT wire_y_pipeff_2_w_q_range1769w(0);
	wire_y_pipeff_2_w_lg_w_q_range1775w1777w(0) <= NOT wire_y_pipeff_2_w_q_range1775w(0);
	wire_y_pipeff_2_w_lg_w_q_range1781w1783w(0) <= NOT wire_y_pipeff_2_w_q_range1781w(0);
	wire_y_pipeff_2_w_lg_w_q_range1787w1789w(0) <= NOT wire_y_pipeff_2_w_q_range1787w(0);
	wire_y_pipeff_2_w_lg_w_q_range1793w1795w(0) <= NOT wire_y_pipeff_2_w_q_range1793w(0);
	wire_y_pipeff_2_w_lg_w_q_range1799w1801w(0) <= NOT wire_y_pipeff_2_w_q_range1799w(0);
	wire_y_pipeff_2_w_lg_w_q_range1805w1807w(0) <= NOT wire_y_pipeff_2_w_q_range1805w(0);
	wire_y_pipeff_2_w_lg_w_q_range1811w1813w(0) <= NOT wire_y_pipeff_2_w_q_range1811w(0);
	wire_y_pipeff_2_w_lg_w_q_range1817w1819w(0) <= NOT wire_y_pipeff_2_w_q_range1817w(0);
	wire_y_pipeff_2_w_lg_w_q_range1823w1825w(0) <= NOT wire_y_pipeff_2_w_q_range1823w(0);
	wire_y_pipeff_2_w_lg_w_q_range1829w1831w(0) <= NOT wire_y_pipeff_2_w_q_range1829w(0);
	wire_y_pipeff_2_w_lg_w_q_range1835w1837w(0) <= NOT wire_y_pipeff_2_w_q_range1835w(0);
	wire_y_pipeff_2_w_lg_w_q_range1841w1843w(0) <= NOT wire_y_pipeff_2_w_q_range1841w(0);
	wire_y_pipeff_2_w_lg_w_q_range1847w1849w(0) <= NOT wire_y_pipeff_2_w_q_range1847w(0);
	wire_y_pipeff_2_w_lg_w_q_range1853w1855w(0) <= NOT wire_y_pipeff_2_w_q_range1853w(0);
	wire_y_pipeff_2_w_lg_w_q_range1859w1861w(0) <= NOT wire_y_pipeff_2_w_q_range1859w(0);
	wire_y_pipeff_2_w_lg_w_q_range1865w1867w(0) <= NOT wire_y_pipeff_2_w_q_range1865w(0);
	wire_y_pipeff_2_w_lg_w_q_range1871w1873w(0) <= NOT wire_y_pipeff_2_w_q_range1871w(0);
	wire_y_pipeff_2_w_lg_w_q_range1877w1879w(0) <= NOT wire_y_pipeff_2_w_q_range1877w(0);
	wire_y_pipeff_2_w_lg_w_q_range1716w1718w(0) <= NOT wire_y_pipeff_2_w_q_range1716w(0);
	wire_y_pipeff_2_w_lg_w_q_range1883w1885w(0) <= NOT wire_y_pipeff_2_w_q_range1883w(0);
	wire_y_pipeff_2_w_lg_w_q_range1889w1891w(0) <= NOT wire_y_pipeff_2_w_q_range1889w(0);
	wire_y_pipeff_2_w_lg_w_q_range1895w1897w(0) <= NOT wire_y_pipeff_2_w_q_range1895w(0);
	wire_y_pipeff_2_w_lg_w_q_range1697w1699w(0) <= NOT wire_y_pipeff_2_w_q_range1697w(0);
	wire_y_pipeff_2_w_lg_w_q_range1721w1723w(0) <= NOT wire_y_pipeff_2_w_q_range1721w(0);
	wire_y_pipeff_2_w_lg_w_q_range1727w1729w(0) <= NOT wire_y_pipeff_2_w_q_range1727w(0);
	wire_y_pipeff_2_w_lg_w_q_range1733w1735w(0) <= NOT wire_y_pipeff_2_w_q_range1733w(0);
	wire_y_pipeff_2_w_lg_w_q_range1739w1741w(0) <= NOT wire_y_pipeff_2_w_q_range1739w(0);
	wire_y_pipeff_2_w_lg_w_q_range1745w1747w(0) <= NOT wire_y_pipeff_2_w_q_range1745w(0);
	wire_y_pipeff_2_w_lg_w_q_range1751w1753w(0) <= NOT wire_y_pipeff_2_w_q_range1751w(0);
	wire_y_pipeff_2_w_lg_w_q_range1757w1759w(0) <= NOT wire_y_pipeff_2_w_q_range1757w(0);
	wire_y_pipeff_2_w_q_range1763w(0) <= y_pipeff_2(10);
	wire_y_pipeff_2_w_q_range1769w(0) <= y_pipeff_2(11);
	wire_y_pipeff_2_w_q_range1775w(0) <= y_pipeff_2(12);
	wire_y_pipeff_2_w_q_range1781w(0) <= y_pipeff_2(13);
	wire_y_pipeff_2_w_q_range1787w(0) <= y_pipeff_2(14);
	wire_y_pipeff_2_w_q_range1793w(0) <= y_pipeff_2(15);
	wire_y_pipeff_2_w_q_range1799w(0) <= y_pipeff_2(16);
	wire_y_pipeff_2_w_q_range1805w(0) <= y_pipeff_2(17);
	wire_y_pipeff_2_w_q_range1811w(0) <= y_pipeff_2(18);
	wire_y_pipeff_2_w_q_range1817w(0) <= y_pipeff_2(19);
	wire_y_pipeff_2_w_q_range1823w(0) <= y_pipeff_2(20);
	wire_y_pipeff_2_w_q_range1829w(0) <= y_pipeff_2(21);
	wire_y_pipeff_2_w_q_range1835w(0) <= y_pipeff_2(22);
	wire_y_pipeff_2_w_q_range1841w(0) <= y_pipeff_2(23);
	wire_y_pipeff_2_w_q_range1847w(0) <= y_pipeff_2(24);
	wire_y_pipeff_2_w_q_range1853w(0) <= y_pipeff_2(25);
	wire_y_pipeff_2_w_q_range1859w(0) <= y_pipeff_2(26);
	wire_y_pipeff_2_w_q_range1865w(0) <= y_pipeff_2(27);
	wire_y_pipeff_2_w_q_range1871w(0) <= y_pipeff_2(28);
	wire_y_pipeff_2_w_q_range1877w(0) <= y_pipeff_2(29);
	wire_y_pipeff_2_w_q_range1716w(0) <= y_pipeff_2(2);
	wire_y_pipeff_2_w_q_range1883w(0) <= y_pipeff_2(30);
	wire_y_pipeff_2_w_q_range1889w(0) <= y_pipeff_2(31);
	wire_y_pipeff_2_w_q_range1895w(0) <= y_pipeff_2(32);
	wire_y_pipeff_2_w_q_range1697w(0) <= y_pipeff_2(33);
	wire_y_pipeff_2_w_q_range1721w(0) <= y_pipeff_2(3);
	wire_y_pipeff_2_w_q_range1727w(0) <= y_pipeff_2(4);
	wire_y_pipeff_2_w_q_range1733w(0) <= y_pipeff_2(5);
	wire_y_pipeff_2_w_q_range1739w(0) <= y_pipeff_2(6);
	wire_y_pipeff_2_w_q_range1745w(0) <= y_pipeff_2(7);
	wire_y_pipeff_2_w_q_range1751w(0) <= y_pipeff_2(8);
	wire_y_pipeff_2_w_q_range1757w(0) <= y_pipeff_2(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_3 <= y_pipenode_3_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_3_w_lg_w_q_range2608w2610w(0) <= NOT wire_y_pipeff_3_w_q_range2608w(0);
	wire_y_pipeff_3_w_lg_w_q_range2614w2616w(0) <= NOT wire_y_pipeff_3_w_q_range2614w(0);
	wire_y_pipeff_3_w_lg_w_q_range2620w2622w(0) <= NOT wire_y_pipeff_3_w_q_range2620w(0);
	wire_y_pipeff_3_w_lg_w_q_range2626w2628w(0) <= NOT wire_y_pipeff_3_w_q_range2626w(0);
	wire_y_pipeff_3_w_lg_w_q_range2632w2634w(0) <= NOT wire_y_pipeff_3_w_q_range2632w(0);
	wire_y_pipeff_3_w_lg_w_q_range2638w2640w(0) <= NOT wire_y_pipeff_3_w_q_range2638w(0);
	wire_y_pipeff_3_w_lg_w_q_range2644w2646w(0) <= NOT wire_y_pipeff_3_w_q_range2644w(0);
	wire_y_pipeff_3_w_lg_w_q_range2650w2652w(0) <= NOT wire_y_pipeff_3_w_q_range2650w(0);
	wire_y_pipeff_3_w_lg_w_q_range2656w2658w(0) <= NOT wire_y_pipeff_3_w_q_range2656w(0);
	wire_y_pipeff_3_w_lg_w_q_range2662w2664w(0) <= NOT wire_y_pipeff_3_w_q_range2662w(0);
	wire_y_pipeff_3_w_lg_w_q_range2668w2670w(0) <= NOT wire_y_pipeff_3_w_q_range2668w(0);
	wire_y_pipeff_3_w_lg_w_q_range2674w2676w(0) <= NOT wire_y_pipeff_3_w_q_range2674w(0);
	wire_y_pipeff_3_w_lg_w_q_range2680w2682w(0) <= NOT wire_y_pipeff_3_w_q_range2680w(0);
	wire_y_pipeff_3_w_lg_w_q_range2686w2688w(0) <= NOT wire_y_pipeff_3_w_q_range2686w(0);
	wire_y_pipeff_3_w_lg_w_q_range2692w2694w(0) <= NOT wire_y_pipeff_3_w_q_range2692w(0);
	wire_y_pipeff_3_w_lg_w_q_range2698w2700w(0) <= NOT wire_y_pipeff_3_w_q_range2698w(0);
	wire_y_pipeff_3_w_lg_w_q_range2704w2706w(0) <= NOT wire_y_pipeff_3_w_q_range2704w(0);
	wire_y_pipeff_3_w_lg_w_q_range2710w2712w(0) <= NOT wire_y_pipeff_3_w_q_range2710w(0);
	wire_y_pipeff_3_w_lg_w_q_range2716w2718w(0) <= NOT wire_y_pipeff_3_w_q_range2716w(0);
	wire_y_pipeff_3_w_lg_w_q_range2722w2724w(0) <= NOT wire_y_pipeff_3_w_q_range2722w(0);
	wire_y_pipeff_3_w_lg_w_q_range2728w2730w(0) <= NOT wire_y_pipeff_3_w_q_range2728w(0);
	wire_y_pipeff_3_w_lg_w_q_range2734w2736w(0) <= NOT wire_y_pipeff_3_w_q_range2734w(0);
	wire_y_pipeff_3_w_lg_w_q_range2740w2742w(0) <= NOT wire_y_pipeff_3_w_q_range2740w(0);
	wire_y_pipeff_3_w_lg_w_q_range2544w2546w(0) <= NOT wire_y_pipeff_3_w_q_range2544w(0);
	wire_y_pipeff_3_w_lg_w_q_range2567w2569w(0) <= NOT wire_y_pipeff_3_w_q_range2567w(0);
	wire_y_pipeff_3_w_lg_w_q_range2572w2574w(0) <= NOT wire_y_pipeff_3_w_q_range2572w(0);
	wire_y_pipeff_3_w_lg_w_q_range2578w2580w(0) <= NOT wire_y_pipeff_3_w_q_range2578w(0);
	wire_y_pipeff_3_w_lg_w_q_range2584w2586w(0) <= NOT wire_y_pipeff_3_w_q_range2584w(0);
	wire_y_pipeff_3_w_lg_w_q_range2590w2592w(0) <= NOT wire_y_pipeff_3_w_q_range2590w(0);
	wire_y_pipeff_3_w_lg_w_q_range2596w2598w(0) <= NOT wire_y_pipeff_3_w_q_range2596w(0);
	wire_y_pipeff_3_w_lg_w_q_range2602w2604w(0) <= NOT wire_y_pipeff_3_w_q_range2602w(0);
	wire_y_pipeff_3_w_q_range2608w(0) <= y_pipeff_3(10);
	wire_y_pipeff_3_w_q_range2614w(0) <= y_pipeff_3(11);
	wire_y_pipeff_3_w_q_range2620w(0) <= y_pipeff_3(12);
	wire_y_pipeff_3_w_q_range2626w(0) <= y_pipeff_3(13);
	wire_y_pipeff_3_w_q_range2632w(0) <= y_pipeff_3(14);
	wire_y_pipeff_3_w_q_range2638w(0) <= y_pipeff_3(15);
	wire_y_pipeff_3_w_q_range2644w(0) <= y_pipeff_3(16);
	wire_y_pipeff_3_w_q_range2650w(0) <= y_pipeff_3(17);
	wire_y_pipeff_3_w_q_range2656w(0) <= y_pipeff_3(18);
	wire_y_pipeff_3_w_q_range2662w(0) <= y_pipeff_3(19);
	wire_y_pipeff_3_w_q_range2668w(0) <= y_pipeff_3(20);
	wire_y_pipeff_3_w_q_range2674w(0) <= y_pipeff_3(21);
	wire_y_pipeff_3_w_q_range2680w(0) <= y_pipeff_3(22);
	wire_y_pipeff_3_w_q_range2686w(0) <= y_pipeff_3(23);
	wire_y_pipeff_3_w_q_range2692w(0) <= y_pipeff_3(24);
	wire_y_pipeff_3_w_q_range2698w(0) <= y_pipeff_3(25);
	wire_y_pipeff_3_w_q_range2704w(0) <= y_pipeff_3(26);
	wire_y_pipeff_3_w_q_range2710w(0) <= y_pipeff_3(27);
	wire_y_pipeff_3_w_q_range2716w(0) <= y_pipeff_3(28);
	wire_y_pipeff_3_w_q_range2722w(0) <= y_pipeff_3(29);
	wire_y_pipeff_3_w_q_range2728w(0) <= y_pipeff_3(30);
	wire_y_pipeff_3_w_q_range2734w(0) <= y_pipeff_3(31);
	wire_y_pipeff_3_w_q_range2740w(0) <= y_pipeff_3(32);
	wire_y_pipeff_3_w_q_range2544w(0) <= y_pipeff_3(33);
	wire_y_pipeff_3_w_q_range2567w(0) <= y_pipeff_3(3);
	wire_y_pipeff_3_w_q_range2572w(0) <= y_pipeff_3(4);
	wire_y_pipeff_3_w_q_range2578w(0) <= y_pipeff_3(5);
	wire_y_pipeff_3_w_q_range2584w(0) <= y_pipeff_3(6);
	wire_y_pipeff_3_w_q_range2590w(0) <= y_pipeff_3(7);
	wire_y_pipeff_3_w_q_range2596w(0) <= y_pipeff_3(8);
	wire_y_pipeff_3_w_q_range2602w(0) <= y_pipeff_3(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_4 <= y_pipenode_4_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_4_w_lg_w_q_range3448w3450w(0) <= NOT wire_y_pipeff_4_w_q_range3448w(0);
	wire_y_pipeff_4_w_lg_w_q_range3454w3456w(0) <= NOT wire_y_pipeff_4_w_q_range3454w(0);
	wire_y_pipeff_4_w_lg_w_q_range3460w3462w(0) <= NOT wire_y_pipeff_4_w_q_range3460w(0);
	wire_y_pipeff_4_w_lg_w_q_range3466w3468w(0) <= NOT wire_y_pipeff_4_w_q_range3466w(0);
	wire_y_pipeff_4_w_lg_w_q_range3472w3474w(0) <= NOT wire_y_pipeff_4_w_q_range3472w(0);
	wire_y_pipeff_4_w_lg_w_q_range3478w3480w(0) <= NOT wire_y_pipeff_4_w_q_range3478w(0);
	wire_y_pipeff_4_w_lg_w_q_range3484w3486w(0) <= NOT wire_y_pipeff_4_w_q_range3484w(0);
	wire_y_pipeff_4_w_lg_w_q_range3490w3492w(0) <= NOT wire_y_pipeff_4_w_q_range3490w(0);
	wire_y_pipeff_4_w_lg_w_q_range3496w3498w(0) <= NOT wire_y_pipeff_4_w_q_range3496w(0);
	wire_y_pipeff_4_w_lg_w_q_range3502w3504w(0) <= NOT wire_y_pipeff_4_w_q_range3502w(0);
	wire_y_pipeff_4_w_lg_w_q_range3508w3510w(0) <= NOT wire_y_pipeff_4_w_q_range3508w(0);
	wire_y_pipeff_4_w_lg_w_q_range3514w3516w(0) <= NOT wire_y_pipeff_4_w_q_range3514w(0);
	wire_y_pipeff_4_w_lg_w_q_range3520w3522w(0) <= NOT wire_y_pipeff_4_w_q_range3520w(0);
	wire_y_pipeff_4_w_lg_w_q_range3526w3528w(0) <= NOT wire_y_pipeff_4_w_q_range3526w(0);
	wire_y_pipeff_4_w_lg_w_q_range3532w3534w(0) <= NOT wire_y_pipeff_4_w_q_range3532w(0);
	wire_y_pipeff_4_w_lg_w_q_range3538w3540w(0) <= NOT wire_y_pipeff_4_w_q_range3538w(0);
	wire_y_pipeff_4_w_lg_w_q_range3544w3546w(0) <= NOT wire_y_pipeff_4_w_q_range3544w(0);
	wire_y_pipeff_4_w_lg_w_q_range3550w3552w(0) <= NOT wire_y_pipeff_4_w_q_range3550w(0);
	wire_y_pipeff_4_w_lg_w_q_range3556w3558w(0) <= NOT wire_y_pipeff_4_w_q_range3556w(0);
	wire_y_pipeff_4_w_lg_w_q_range3562w3564w(0) <= NOT wire_y_pipeff_4_w_q_range3562w(0);
	wire_y_pipeff_4_w_lg_w_q_range3568w3570w(0) <= NOT wire_y_pipeff_4_w_q_range3568w(0);
	wire_y_pipeff_4_w_lg_w_q_range3574w3576w(0) <= NOT wire_y_pipeff_4_w_q_range3574w(0);
	wire_y_pipeff_4_w_lg_w_q_range3580w3582w(0) <= NOT wire_y_pipeff_4_w_q_range3580w(0);
	wire_y_pipeff_4_w_lg_w_q_range3386w3388w(0) <= NOT wire_y_pipeff_4_w_q_range3386w(0);
	wire_y_pipeff_4_w_lg_w_q_range3413w3415w(0) <= NOT wire_y_pipeff_4_w_q_range3413w(0);
	wire_y_pipeff_4_w_lg_w_q_range3418w3420w(0) <= NOT wire_y_pipeff_4_w_q_range3418w(0);
	wire_y_pipeff_4_w_lg_w_q_range3424w3426w(0) <= NOT wire_y_pipeff_4_w_q_range3424w(0);
	wire_y_pipeff_4_w_lg_w_q_range3430w3432w(0) <= NOT wire_y_pipeff_4_w_q_range3430w(0);
	wire_y_pipeff_4_w_lg_w_q_range3436w3438w(0) <= NOT wire_y_pipeff_4_w_q_range3436w(0);
	wire_y_pipeff_4_w_lg_w_q_range3442w3444w(0) <= NOT wire_y_pipeff_4_w_q_range3442w(0);
	wire_y_pipeff_4_w_q_range3448w(0) <= y_pipeff_4(10);
	wire_y_pipeff_4_w_q_range3454w(0) <= y_pipeff_4(11);
	wire_y_pipeff_4_w_q_range3460w(0) <= y_pipeff_4(12);
	wire_y_pipeff_4_w_q_range3466w(0) <= y_pipeff_4(13);
	wire_y_pipeff_4_w_q_range3472w(0) <= y_pipeff_4(14);
	wire_y_pipeff_4_w_q_range3478w(0) <= y_pipeff_4(15);
	wire_y_pipeff_4_w_q_range3484w(0) <= y_pipeff_4(16);
	wire_y_pipeff_4_w_q_range3490w(0) <= y_pipeff_4(17);
	wire_y_pipeff_4_w_q_range3496w(0) <= y_pipeff_4(18);
	wire_y_pipeff_4_w_q_range3502w(0) <= y_pipeff_4(19);
	wire_y_pipeff_4_w_q_range3508w(0) <= y_pipeff_4(20);
	wire_y_pipeff_4_w_q_range3514w(0) <= y_pipeff_4(21);
	wire_y_pipeff_4_w_q_range3520w(0) <= y_pipeff_4(22);
	wire_y_pipeff_4_w_q_range3526w(0) <= y_pipeff_4(23);
	wire_y_pipeff_4_w_q_range3532w(0) <= y_pipeff_4(24);
	wire_y_pipeff_4_w_q_range3538w(0) <= y_pipeff_4(25);
	wire_y_pipeff_4_w_q_range3544w(0) <= y_pipeff_4(26);
	wire_y_pipeff_4_w_q_range3550w(0) <= y_pipeff_4(27);
	wire_y_pipeff_4_w_q_range3556w(0) <= y_pipeff_4(28);
	wire_y_pipeff_4_w_q_range3562w(0) <= y_pipeff_4(29);
	wire_y_pipeff_4_w_q_range3568w(0) <= y_pipeff_4(30);
	wire_y_pipeff_4_w_q_range3574w(0) <= y_pipeff_4(31);
	wire_y_pipeff_4_w_q_range3580w(0) <= y_pipeff_4(32);
	wire_y_pipeff_4_w_q_range3386w(0) <= y_pipeff_4(33);
	wire_y_pipeff_4_w_q_range3413w(0) <= y_pipeff_4(4);
	wire_y_pipeff_4_w_q_range3418w(0) <= y_pipeff_4(5);
	wire_y_pipeff_4_w_q_range3424w(0) <= y_pipeff_4(6);
	wire_y_pipeff_4_w_q_range3430w(0) <= y_pipeff_4(7);
	wire_y_pipeff_4_w_q_range3436w(0) <= y_pipeff_4(8);
	wire_y_pipeff_4_w_q_range3442w(0) <= y_pipeff_4(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_5 <= y_pipenode_5_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_5_w_lg_w_q_range4283w4285w(0) <= NOT wire_y_pipeff_5_w_q_range4283w(0);
	wire_y_pipeff_5_w_lg_w_q_range4289w4291w(0) <= NOT wire_y_pipeff_5_w_q_range4289w(0);
	wire_y_pipeff_5_w_lg_w_q_range4295w4297w(0) <= NOT wire_y_pipeff_5_w_q_range4295w(0);
	wire_y_pipeff_5_w_lg_w_q_range4301w4303w(0) <= NOT wire_y_pipeff_5_w_q_range4301w(0);
	wire_y_pipeff_5_w_lg_w_q_range4307w4309w(0) <= NOT wire_y_pipeff_5_w_q_range4307w(0);
	wire_y_pipeff_5_w_lg_w_q_range4313w4315w(0) <= NOT wire_y_pipeff_5_w_q_range4313w(0);
	wire_y_pipeff_5_w_lg_w_q_range4319w4321w(0) <= NOT wire_y_pipeff_5_w_q_range4319w(0);
	wire_y_pipeff_5_w_lg_w_q_range4325w4327w(0) <= NOT wire_y_pipeff_5_w_q_range4325w(0);
	wire_y_pipeff_5_w_lg_w_q_range4331w4333w(0) <= NOT wire_y_pipeff_5_w_q_range4331w(0);
	wire_y_pipeff_5_w_lg_w_q_range4337w4339w(0) <= NOT wire_y_pipeff_5_w_q_range4337w(0);
	wire_y_pipeff_5_w_lg_w_q_range4343w4345w(0) <= NOT wire_y_pipeff_5_w_q_range4343w(0);
	wire_y_pipeff_5_w_lg_w_q_range4349w4351w(0) <= NOT wire_y_pipeff_5_w_q_range4349w(0);
	wire_y_pipeff_5_w_lg_w_q_range4355w4357w(0) <= NOT wire_y_pipeff_5_w_q_range4355w(0);
	wire_y_pipeff_5_w_lg_w_q_range4361w4363w(0) <= NOT wire_y_pipeff_5_w_q_range4361w(0);
	wire_y_pipeff_5_w_lg_w_q_range4367w4369w(0) <= NOT wire_y_pipeff_5_w_q_range4367w(0);
	wire_y_pipeff_5_w_lg_w_q_range4373w4375w(0) <= NOT wire_y_pipeff_5_w_q_range4373w(0);
	wire_y_pipeff_5_w_lg_w_q_range4379w4381w(0) <= NOT wire_y_pipeff_5_w_q_range4379w(0);
	wire_y_pipeff_5_w_lg_w_q_range4385w4387w(0) <= NOT wire_y_pipeff_5_w_q_range4385w(0);
	wire_y_pipeff_5_w_lg_w_q_range4391w4393w(0) <= NOT wire_y_pipeff_5_w_q_range4391w(0);
	wire_y_pipeff_5_w_lg_w_q_range4397w4399w(0) <= NOT wire_y_pipeff_5_w_q_range4397w(0);
	wire_y_pipeff_5_w_lg_w_q_range4403w4405w(0) <= NOT wire_y_pipeff_5_w_q_range4403w(0);
	wire_y_pipeff_5_w_lg_w_q_range4409w4411w(0) <= NOT wire_y_pipeff_5_w_q_range4409w(0);
	wire_y_pipeff_5_w_lg_w_q_range4415w4417w(0) <= NOT wire_y_pipeff_5_w_q_range4415w(0);
	wire_y_pipeff_5_w_lg_w_q_range4223w4225w(0) <= NOT wire_y_pipeff_5_w_q_range4223w(0);
	wire_y_pipeff_5_w_lg_w_q_range4254w4256w(0) <= NOT wire_y_pipeff_5_w_q_range4254w(0);
	wire_y_pipeff_5_w_lg_w_q_range4259w4261w(0) <= NOT wire_y_pipeff_5_w_q_range4259w(0);
	wire_y_pipeff_5_w_lg_w_q_range4265w4267w(0) <= NOT wire_y_pipeff_5_w_q_range4265w(0);
	wire_y_pipeff_5_w_lg_w_q_range4271w4273w(0) <= NOT wire_y_pipeff_5_w_q_range4271w(0);
	wire_y_pipeff_5_w_lg_w_q_range4277w4279w(0) <= NOT wire_y_pipeff_5_w_q_range4277w(0);
	wire_y_pipeff_5_w_q_range4283w(0) <= y_pipeff_5(10);
	wire_y_pipeff_5_w_q_range4289w(0) <= y_pipeff_5(11);
	wire_y_pipeff_5_w_q_range4295w(0) <= y_pipeff_5(12);
	wire_y_pipeff_5_w_q_range4301w(0) <= y_pipeff_5(13);
	wire_y_pipeff_5_w_q_range4307w(0) <= y_pipeff_5(14);
	wire_y_pipeff_5_w_q_range4313w(0) <= y_pipeff_5(15);
	wire_y_pipeff_5_w_q_range4319w(0) <= y_pipeff_5(16);
	wire_y_pipeff_5_w_q_range4325w(0) <= y_pipeff_5(17);
	wire_y_pipeff_5_w_q_range4331w(0) <= y_pipeff_5(18);
	wire_y_pipeff_5_w_q_range4337w(0) <= y_pipeff_5(19);
	wire_y_pipeff_5_w_q_range4343w(0) <= y_pipeff_5(20);
	wire_y_pipeff_5_w_q_range4349w(0) <= y_pipeff_5(21);
	wire_y_pipeff_5_w_q_range4355w(0) <= y_pipeff_5(22);
	wire_y_pipeff_5_w_q_range4361w(0) <= y_pipeff_5(23);
	wire_y_pipeff_5_w_q_range4367w(0) <= y_pipeff_5(24);
	wire_y_pipeff_5_w_q_range4373w(0) <= y_pipeff_5(25);
	wire_y_pipeff_5_w_q_range4379w(0) <= y_pipeff_5(26);
	wire_y_pipeff_5_w_q_range4385w(0) <= y_pipeff_5(27);
	wire_y_pipeff_5_w_q_range4391w(0) <= y_pipeff_5(28);
	wire_y_pipeff_5_w_q_range4397w(0) <= y_pipeff_5(29);
	wire_y_pipeff_5_w_q_range4403w(0) <= y_pipeff_5(30);
	wire_y_pipeff_5_w_q_range4409w(0) <= y_pipeff_5(31);
	wire_y_pipeff_5_w_q_range4415w(0) <= y_pipeff_5(32);
	wire_y_pipeff_5_w_q_range4223w(0) <= y_pipeff_5(33);
	wire_y_pipeff_5_w_q_range4254w(0) <= y_pipeff_5(5);
	wire_y_pipeff_5_w_q_range4259w(0) <= y_pipeff_5(6);
	wire_y_pipeff_5_w_q_range4265w(0) <= y_pipeff_5(7);
	wire_y_pipeff_5_w_q_range4271w(0) <= y_pipeff_5(8);
	wire_y_pipeff_5_w_q_range4277w(0) <= y_pipeff_5(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_6 <= y_pipenode_6_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_6_w_lg_w_q_range5113w5115w(0) <= NOT wire_y_pipeff_6_w_q_range5113w(0);
	wire_y_pipeff_6_w_lg_w_q_range5119w5121w(0) <= NOT wire_y_pipeff_6_w_q_range5119w(0);
	wire_y_pipeff_6_w_lg_w_q_range5125w5127w(0) <= NOT wire_y_pipeff_6_w_q_range5125w(0);
	wire_y_pipeff_6_w_lg_w_q_range5131w5133w(0) <= NOT wire_y_pipeff_6_w_q_range5131w(0);
	wire_y_pipeff_6_w_lg_w_q_range5137w5139w(0) <= NOT wire_y_pipeff_6_w_q_range5137w(0);
	wire_y_pipeff_6_w_lg_w_q_range5143w5145w(0) <= NOT wire_y_pipeff_6_w_q_range5143w(0);
	wire_y_pipeff_6_w_lg_w_q_range5149w5151w(0) <= NOT wire_y_pipeff_6_w_q_range5149w(0);
	wire_y_pipeff_6_w_lg_w_q_range5155w5157w(0) <= NOT wire_y_pipeff_6_w_q_range5155w(0);
	wire_y_pipeff_6_w_lg_w_q_range5161w5163w(0) <= NOT wire_y_pipeff_6_w_q_range5161w(0);
	wire_y_pipeff_6_w_lg_w_q_range5167w5169w(0) <= NOT wire_y_pipeff_6_w_q_range5167w(0);
	wire_y_pipeff_6_w_lg_w_q_range5173w5175w(0) <= NOT wire_y_pipeff_6_w_q_range5173w(0);
	wire_y_pipeff_6_w_lg_w_q_range5179w5181w(0) <= NOT wire_y_pipeff_6_w_q_range5179w(0);
	wire_y_pipeff_6_w_lg_w_q_range5185w5187w(0) <= NOT wire_y_pipeff_6_w_q_range5185w(0);
	wire_y_pipeff_6_w_lg_w_q_range5191w5193w(0) <= NOT wire_y_pipeff_6_w_q_range5191w(0);
	wire_y_pipeff_6_w_lg_w_q_range5197w5199w(0) <= NOT wire_y_pipeff_6_w_q_range5197w(0);
	wire_y_pipeff_6_w_lg_w_q_range5203w5205w(0) <= NOT wire_y_pipeff_6_w_q_range5203w(0);
	wire_y_pipeff_6_w_lg_w_q_range5209w5211w(0) <= NOT wire_y_pipeff_6_w_q_range5209w(0);
	wire_y_pipeff_6_w_lg_w_q_range5215w5217w(0) <= NOT wire_y_pipeff_6_w_q_range5215w(0);
	wire_y_pipeff_6_w_lg_w_q_range5221w5223w(0) <= NOT wire_y_pipeff_6_w_q_range5221w(0);
	wire_y_pipeff_6_w_lg_w_q_range5227w5229w(0) <= NOT wire_y_pipeff_6_w_q_range5227w(0);
	wire_y_pipeff_6_w_lg_w_q_range5233w5235w(0) <= NOT wire_y_pipeff_6_w_q_range5233w(0);
	wire_y_pipeff_6_w_lg_w_q_range5239w5241w(0) <= NOT wire_y_pipeff_6_w_q_range5239w(0);
	wire_y_pipeff_6_w_lg_w_q_range5245w5247w(0) <= NOT wire_y_pipeff_6_w_q_range5245w(0);
	wire_y_pipeff_6_w_lg_w_q_range5055w5057w(0) <= NOT wire_y_pipeff_6_w_q_range5055w(0);
	wire_y_pipeff_6_w_lg_w_q_range5090w5092w(0) <= NOT wire_y_pipeff_6_w_q_range5090w(0);
	wire_y_pipeff_6_w_lg_w_q_range5095w5097w(0) <= NOT wire_y_pipeff_6_w_q_range5095w(0);
	wire_y_pipeff_6_w_lg_w_q_range5101w5103w(0) <= NOT wire_y_pipeff_6_w_q_range5101w(0);
	wire_y_pipeff_6_w_lg_w_q_range5107w5109w(0) <= NOT wire_y_pipeff_6_w_q_range5107w(0);
	wire_y_pipeff_6_w_q_range5113w(0) <= y_pipeff_6(10);
	wire_y_pipeff_6_w_q_range5119w(0) <= y_pipeff_6(11);
	wire_y_pipeff_6_w_q_range5125w(0) <= y_pipeff_6(12);
	wire_y_pipeff_6_w_q_range5131w(0) <= y_pipeff_6(13);
	wire_y_pipeff_6_w_q_range5137w(0) <= y_pipeff_6(14);
	wire_y_pipeff_6_w_q_range5143w(0) <= y_pipeff_6(15);
	wire_y_pipeff_6_w_q_range5149w(0) <= y_pipeff_6(16);
	wire_y_pipeff_6_w_q_range5155w(0) <= y_pipeff_6(17);
	wire_y_pipeff_6_w_q_range5161w(0) <= y_pipeff_6(18);
	wire_y_pipeff_6_w_q_range5167w(0) <= y_pipeff_6(19);
	wire_y_pipeff_6_w_q_range5173w(0) <= y_pipeff_6(20);
	wire_y_pipeff_6_w_q_range5179w(0) <= y_pipeff_6(21);
	wire_y_pipeff_6_w_q_range5185w(0) <= y_pipeff_6(22);
	wire_y_pipeff_6_w_q_range5191w(0) <= y_pipeff_6(23);
	wire_y_pipeff_6_w_q_range5197w(0) <= y_pipeff_6(24);
	wire_y_pipeff_6_w_q_range5203w(0) <= y_pipeff_6(25);
	wire_y_pipeff_6_w_q_range5209w(0) <= y_pipeff_6(26);
	wire_y_pipeff_6_w_q_range5215w(0) <= y_pipeff_6(27);
	wire_y_pipeff_6_w_q_range5221w(0) <= y_pipeff_6(28);
	wire_y_pipeff_6_w_q_range5227w(0) <= y_pipeff_6(29);
	wire_y_pipeff_6_w_q_range5233w(0) <= y_pipeff_6(30);
	wire_y_pipeff_6_w_q_range5239w(0) <= y_pipeff_6(31);
	wire_y_pipeff_6_w_q_range5245w(0) <= y_pipeff_6(32);
	wire_y_pipeff_6_w_q_range5055w(0) <= y_pipeff_6(33);
	wire_y_pipeff_6_w_q_range5090w(0) <= y_pipeff_6(6);
	wire_y_pipeff_6_w_q_range5095w(0) <= y_pipeff_6(7);
	wire_y_pipeff_6_w_q_range5101w(0) <= y_pipeff_6(8);
	wire_y_pipeff_6_w_q_range5107w(0) <= y_pipeff_6(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_7 <= y_pipenode_7_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_7_w_lg_w_q_range5938w5940w(0) <= NOT wire_y_pipeff_7_w_q_range5938w(0);
	wire_y_pipeff_7_w_lg_w_q_range5944w5946w(0) <= NOT wire_y_pipeff_7_w_q_range5944w(0);
	wire_y_pipeff_7_w_lg_w_q_range5950w5952w(0) <= NOT wire_y_pipeff_7_w_q_range5950w(0);
	wire_y_pipeff_7_w_lg_w_q_range5956w5958w(0) <= NOT wire_y_pipeff_7_w_q_range5956w(0);
	wire_y_pipeff_7_w_lg_w_q_range5962w5964w(0) <= NOT wire_y_pipeff_7_w_q_range5962w(0);
	wire_y_pipeff_7_w_lg_w_q_range5968w5970w(0) <= NOT wire_y_pipeff_7_w_q_range5968w(0);
	wire_y_pipeff_7_w_lg_w_q_range5974w5976w(0) <= NOT wire_y_pipeff_7_w_q_range5974w(0);
	wire_y_pipeff_7_w_lg_w_q_range5980w5982w(0) <= NOT wire_y_pipeff_7_w_q_range5980w(0);
	wire_y_pipeff_7_w_lg_w_q_range5986w5988w(0) <= NOT wire_y_pipeff_7_w_q_range5986w(0);
	wire_y_pipeff_7_w_lg_w_q_range5992w5994w(0) <= NOT wire_y_pipeff_7_w_q_range5992w(0);
	wire_y_pipeff_7_w_lg_w_q_range5998w6000w(0) <= NOT wire_y_pipeff_7_w_q_range5998w(0);
	wire_y_pipeff_7_w_lg_w_q_range6004w6006w(0) <= NOT wire_y_pipeff_7_w_q_range6004w(0);
	wire_y_pipeff_7_w_lg_w_q_range6010w6012w(0) <= NOT wire_y_pipeff_7_w_q_range6010w(0);
	wire_y_pipeff_7_w_lg_w_q_range6016w6018w(0) <= NOT wire_y_pipeff_7_w_q_range6016w(0);
	wire_y_pipeff_7_w_lg_w_q_range6022w6024w(0) <= NOT wire_y_pipeff_7_w_q_range6022w(0);
	wire_y_pipeff_7_w_lg_w_q_range6028w6030w(0) <= NOT wire_y_pipeff_7_w_q_range6028w(0);
	wire_y_pipeff_7_w_lg_w_q_range6034w6036w(0) <= NOT wire_y_pipeff_7_w_q_range6034w(0);
	wire_y_pipeff_7_w_lg_w_q_range6040w6042w(0) <= NOT wire_y_pipeff_7_w_q_range6040w(0);
	wire_y_pipeff_7_w_lg_w_q_range6046w6048w(0) <= NOT wire_y_pipeff_7_w_q_range6046w(0);
	wire_y_pipeff_7_w_lg_w_q_range6052w6054w(0) <= NOT wire_y_pipeff_7_w_q_range6052w(0);
	wire_y_pipeff_7_w_lg_w_q_range6058w6060w(0) <= NOT wire_y_pipeff_7_w_q_range6058w(0);
	wire_y_pipeff_7_w_lg_w_q_range6064w6066w(0) <= NOT wire_y_pipeff_7_w_q_range6064w(0);
	wire_y_pipeff_7_w_lg_w_q_range6070w6072w(0) <= NOT wire_y_pipeff_7_w_q_range6070w(0);
	wire_y_pipeff_7_w_lg_w_q_range5882w5884w(0) <= NOT wire_y_pipeff_7_w_q_range5882w(0);
	wire_y_pipeff_7_w_lg_w_q_range5921w5923w(0) <= NOT wire_y_pipeff_7_w_q_range5921w(0);
	wire_y_pipeff_7_w_lg_w_q_range5926w5928w(0) <= NOT wire_y_pipeff_7_w_q_range5926w(0);
	wire_y_pipeff_7_w_lg_w_q_range5932w5934w(0) <= NOT wire_y_pipeff_7_w_q_range5932w(0);
	wire_y_pipeff_7_w_q_range5938w(0) <= y_pipeff_7(10);
	wire_y_pipeff_7_w_q_range5944w(0) <= y_pipeff_7(11);
	wire_y_pipeff_7_w_q_range5950w(0) <= y_pipeff_7(12);
	wire_y_pipeff_7_w_q_range5956w(0) <= y_pipeff_7(13);
	wire_y_pipeff_7_w_q_range5962w(0) <= y_pipeff_7(14);
	wire_y_pipeff_7_w_q_range5968w(0) <= y_pipeff_7(15);
	wire_y_pipeff_7_w_q_range5974w(0) <= y_pipeff_7(16);
	wire_y_pipeff_7_w_q_range5980w(0) <= y_pipeff_7(17);
	wire_y_pipeff_7_w_q_range5986w(0) <= y_pipeff_7(18);
	wire_y_pipeff_7_w_q_range5992w(0) <= y_pipeff_7(19);
	wire_y_pipeff_7_w_q_range5998w(0) <= y_pipeff_7(20);
	wire_y_pipeff_7_w_q_range6004w(0) <= y_pipeff_7(21);
	wire_y_pipeff_7_w_q_range6010w(0) <= y_pipeff_7(22);
	wire_y_pipeff_7_w_q_range6016w(0) <= y_pipeff_7(23);
	wire_y_pipeff_7_w_q_range6022w(0) <= y_pipeff_7(24);
	wire_y_pipeff_7_w_q_range6028w(0) <= y_pipeff_7(25);
	wire_y_pipeff_7_w_q_range6034w(0) <= y_pipeff_7(26);
	wire_y_pipeff_7_w_q_range6040w(0) <= y_pipeff_7(27);
	wire_y_pipeff_7_w_q_range6046w(0) <= y_pipeff_7(28);
	wire_y_pipeff_7_w_q_range6052w(0) <= y_pipeff_7(29);
	wire_y_pipeff_7_w_q_range6058w(0) <= y_pipeff_7(30);
	wire_y_pipeff_7_w_q_range6064w(0) <= y_pipeff_7(31);
	wire_y_pipeff_7_w_q_range6070w(0) <= y_pipeff_7(32);
	wire_y_pipeff_7_w_q_range5882w(0) <= y_pipeff_7(33);
	wire_y_pipeff_7_w_q_range5921w(0) <= y_pipeff_7(7);
	wire_y_pipeff_7_w_q_range5926w(0) <= y_pipeff_7(8);
	wire_y_pipeff_7_w_q_range5932w(0) <= y_pipeff_7(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_8 <= y_pipenode_8_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_8_w_lg_w_q_range6758w6760w(0) <= NOT wire_y_pipeff_8_w_q_range6758w(0);
	wire_y_pipeff_8_w_lg_w_q_range6764w6766w(0) <= NOT wire_y_pipeff_8_w_q_range6764w(0);
	wire_y_pipeff_8_w_lg_w_q_range6770w6772w(0) <= NOT wire_y_pipeff_8_w_q_range6770w(0);
	wire_y_pipeff_8_w_lg_w_q_range6776w6778w(0) <= NOT wire_y_pipeff_8_w_q_range6776w(0);
	wire_y_pipeff_8_w_lg_w_q_range6782w6784w(0) <= NOT wire_y_pipeff_8_w_q_range6782w(0);
	wire_y_pipeff_8_w_lg_w_q_range6788w6790w(0) <= NOT wire_y_pipeff_8_w_q_range6788w(0);
	wire_y_pipeff_8_w_lg_w_q_range6794w6796w(0) <= NOT wire_y_pipeff_8_w_q_range6794w(0);
	wire_y_pipeff_8_w_lg_w_q_range6800w6802w(0) <= NOT wire_y_pipeff_8_w_q_range6800w(0);
	wire_y_pipeff_8_w_lg_w_q_range6806w6808w(0) <= NOT wire_y_pipeff_8_w_q_range6806w(0);
	wire_y_pipeff_8_w_lg_w_q_range6812w6814w(0) <= NOT wire_y_pipeff_8_w_q_range6812w(0);
	wire_y_pipeff_8_w_lg_w_q_range6818w6820w(0) <= NOT wire_y_pipeff_8_w_q_range6818w(0);
	wire_y_pipeff_8_w_lg_w_q_range6824w6826w(0) <= NOT wire_y_pipeff_8_w_q_range6824w(0);
	wire_y_pipeff_8_w_lg_w_q_range6830w6832w(0) <= NOT wire_y_pipeff_8_w_q_range6830w(0);
	wire_y_pipeff_8_w_lg_w_q_range6836w6838w(0) <= NOT wire_y_pipeff_8_w_q_range6836w(0);
	wire_y_pipeff_8_w_lg_w_q_range6842w6844w(0) <= NOT wire_y_pipeff_8_w_q_range6842w(0);
	wire_y_pipeff_8_w_lg_w_q_range6848w6850w(0) <= NOT wire_y_pipeff_8_w_q_range6848w(0);
	wire_y_pipeff_8_w_lg_w_q_range6854w6856w(0) <= NOT wire_y_pipeff_8_w_q_range6854w(0);
	wire_y_pipeff_8_w_lg_w_q_range6860w6862w(0) <= NOT wire_y_pipeff_8_w_q_range6860w(0);
	wire_y_pipeff_8_w_lg_w_q_range6866w6868w(0) <= NOT wire_y_pipeff_8_w_q_range6866w(0);
	wire_y_pipeff_8_w_lg_w_q_range6872w6874w(0) <= NOT wire_y_pipeff_8_w_q_range6872w(0);
	wire_y_pipeff_8_w_lg_w_q_range6878w6880w(0) <= NOT wire_y_pipeff_8_w_q_range6878w(0);
	wire_y_pipeff_8_w_lg_w_q_range6884w6886w(0) <= NOT wire_y_pipeff_8_w_q_range6884w(0);
	wire_y_pipeff_8_w_lg_w_q_range6890w6892w(0) <= NOT wire_y_pipeff_8_w_q_range6890w(0);
	wire_y_pipeff_8_w_lg_w_q_range6704w6706w(0) <= NOT wire_y_pipeff_8_w_q_range6704w(0);
	wire_y_pipeff_8_w_lg_w_q_range6747w6749w(0) <= NOT wire_y_pipeff_8_w_q_range6747w(0);
	wire_y_pipeff_8_w_lg_w_q_range6752w6754w(0) <= NOT wire_y_pipeff_8_w_q_range6752w(0);
	wire_y_pipeff_8_w_q_range6758w(0) <= y_pipeff_8(10);
	wire_y_pipeff_8_w_q_range6764w(0) <= y_pipeff_8(11);
	wire_y_pipeff_8_w_q_range6770w(0) <= y_pipeff_8(12);
	wire_y_pipeff_8_w_q_range6776w(0) <= y_pipeff_8(13);
	wire_y_pipeff_8_w_q_range6782w(0) <= y_pipeff_8(14);
	wire_y_pipeff_8_w_q_range6788w(0) <= y_pipeff_8(15);
	wire_y_pipeff_8_w_q_range6794w(0) <= y_pipeff_8(16);
	wire_y_pipeff_8_w_q_range6800w(0) <= y_pipeff_8(17);
	wire_y_pipeff_8_w_q_range6806w(0) <= y_pipeff_8(18);
	wire_y_pipeff_8_w_q_range6812w(0) <= y_pipeff_8(19);
	wire_y_pipeff_8_w_q_range6818w(0) <= y_pipeff_8(20);
	wire_y_pipeff_8_w_q_range6824w(0) <= y_pipeff_8(21);
	wire_y_pipeff_8_w_q_range6830w(0) <= y_pipeff_8(22);
	wire_y_pipeff_8_w_q_range6836w(0) <= y_pipeff_8(23);
	wire_y_pipeff_8_w_q_range6842w(0) <= y_pipeff_8(24);
	wire_y_pipeff_8_w_q_range6848w(0) <= y_pipeff_8(25);
	wire_y_pipeff_8_w_q_range6854w(0) <= y_pipeff_8(26);
	wire_y_pipeff_8_w_q_range6860w(0) <= y_pipeff_8(27);
	wire_y_pipeff_8_w_q_range6866w(0) <= y_pipeff_8(28);
	wire_y_pipeff_8_w_q_range6872w(0) <= y_pipeff_8(29);
	wire_y_pipeff_8_w_q_range6878w(0) <= y_pipeff_8(30);
	wire_y_pipeff_8_w_q_range6884w(0) <= y_pipeff_8(31);
	wire_y_pipeff_8_w_q_range6890w(0) <= y_pipeff_8(32);
	wire_y_pipeff_8_w_q_range6704w(0) <= y_pipeff_8(33);
	wire_y_pipeff_8_w_q_range6747w(0) <= y_pipeff_8(8);
	wire_y_pipeff_8_w_q_range6752w(0) <= y_pipeff_8(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_9 <= y_pipenode_9_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_9_w_lg_w_q_range7573w7575w(0) <= NOT wire_y_pipeff_9_w_q_range7573w(0);
	wire_y_pipeff_9_w_lg_w_q_range7579w7581w(0) <= NOT wire_y_pipeff_9_w_q_range7579w(0);
	wire_y_pipeff_9_w_lg_w_q_range7585w7587w(0) <= NOT wire_y_pipeff_9_w_q_range7585w(0);
	wire_y_pipeff_9_w_lg_w_q_range7591w7593w(0) <= NOT wire_y_pipeff_9_w_q_range7591w(0);
	wire_y_pipeff_9_w_lg_w_q_range7597w7599w(0) <= NOT wire_y_pipeff_9_w_q_range7597w(0);
	wire_y_pipeff_9_w_lg_w_q_range7603w7605w(0) <= NOT wire_y_pipeff_9_w_q_range7603w(0);
	wire_y_pipeff_9_w_lg_w_q_range7609w7611w(0) <= NOT wire_y_pipeff_9_w_q_range7609w(0);
	wire_y_pipeff_9_w_lg_w_q_range7615w7617w(0) <= NOT wire_y_pipeff_9_w_q_range7615w(0);
	wire_y_pipeff_9_w_lg_w_q_range7621w7623w(0) <= NOT wire_y_pipeff_9_w_q_range7621w(0);
	wire_y_pipeff_9_w_lg_w_q_range7627w7629w(0) <= NOT wire_y_pipeff_9_w_q_range7627w(0);
	wire_y_pipeff_9_w_lg_w_q_range7633w7635w(0) <= NOT wire_y_pipeff_9_w_q_range7633w(0);
	wire_y_pipeff_9_w_lg_w_q_range7639w7641w(0) <= NOT wire_y_pipeff_9_w_q_range7639w(0);
	wire_y_pipeff_9_w_lg_w_q_range7645w7647w(0) <= NOT wire_y_pipeff_9_w_q_range7645w(0);
	wire_y_pipeff_9_w_lg_w_q_range7651w7653w(0) <= NOT wire_y_pipeff_9_w_q_range7651w(0);
	wire_y_pipeff_9_w_lg_w_q_range7657w7659w(0) <= NOT wire_y_pipeff_9_w_q_range7657w(0);
	wire_y_pipeff_9_w_lg_w_q_range7663w7665w(0) <= NOT wire_y_pipeff_9_w_q_range7663w(0);
	wire_y_pipeff_9_w_lg_w_q_range7669w7671w(0) <= NOT wire_y_pipeff_9_w_q_range7669w(0);
	wire_y_pipeff_9_w_lg_w_q_range7675w7677w(0) <= NOT wire_y_pipeff_9_w_q_range7675w(0);
	wire_y_pipeff_9_w_lg_w_q_range7681w7683w(0) <= NOT wire_y_pipeff_9_w_q_range7681w(0);
	wire_y_pipeff_9_w_lg_w_q_range7687w7689w(0) <= NOT wire_y_pipeff_9_w_q_range7687w(0);
	wire_y_pipeff_9_w_lg_w_q_range7693w7695w(0) <= NOT wire_y_pipeff_9_w_q_range7693w(0);
	wire_y_pipeff_9_w_lg_w_q_range7699w7701w(0) <= NOT wire_y_pipeff_9_w_q_range7699w(0);
	wire_y_pipeff_9_w_lg_w_q_range7705w7707w(0) <= NOT wire_y_pipeff_9_w_q_range7705w(0);
	wire_y_pipeff_9_w_lg_w_q_range7521w7523w(0) <= NOT wire_y_pipeff_9_w_q_range7521w(0);
	wire_y_pipeff_9_w_lg_w_q_range7568w7570w(0) <= NOT wire_y_pipeff_9_w_q_range7568w(0);
	wire_y_pipeff_9_w_q_range7573w(0) <= y_pipeff_9(10);
	wire_y_pipeff_9_w_q_range7579w(0) <= y_pipeff_9(11);
	wire_y_pipeff_9_w_q_range7585w(0) <= y_pipeff_9(12);
	wire_y_pipeff_9_w_q_range7591w(0) <= y_pipeff_9(13);
	wire_y_pipeff_9_w_q_range7597w(0) <= y_pipeff_9(14);
	wire_y_pipeff_9_w_q_range7603w(0) <= y_pipeff_9(15);
	wire_y_pipeff_9_w_q_range7609w(0) <= y_pipeff_9(16);
	wire_y_pipeff_9_w_q_range7615w(0) <= y_pipeff_9(17);
	wire_y_pipeff_9_w_q_range7621w(0) <= y_pipeff_9(18);
	wire_y_pipeff_9_w_q_range7627w(0) <= y_pipeff_9(19);
	wire_y_pipeff_9_w_q_range7633w(0) <= y_pipeff_9(20);
	wire_y_pipeff_9_w_q_range7639w(0) <= y_pipeff_9(21);
	wire_y_pipeff_9_w_q_range7645w(0) <= y_pipeff_9(22);
	wire_y_pipeff_9_w_q_range7651w(0) <= y_pipeff_9(23);
	wire_y_pipeff_9_w_q_range7657w(0) <= y_pipeff_9(24);
	wire_y_pipeff_9_w_q_range7663w(0) <= y_pipeff_9(25);
	wire_y_pipeff_9_w_q_range7669w(0) <= y_pipeff_9(26);
	wire_y_pipeff_9_w_q_range7675w(0) <= y_pipeff_9(27);
	wire_y_pipeff_9_w_q_range7681w(0) <= y_pipeff_9(28);
	wire_y_pipeff_9_w_q_range7687w(0) <= y_pipeff_9(29);
	wire_y_pipeff_9_w_q_range7693w(0) <= y_pipeff_9(30);
	wire_y_pipeff_9_w_q_range7699w(0) <= y_pipeff_9(31);
	wire_y_pipeff_9_w_q_range7705w(0) <= y_pipeff_9(32);
	wire_y_pipeff_9_w_q_range7521w(0) <= y_pipeff_9(33);
	wire_y_pipeff_9_w_q_range7568w(0) <= y_pipeff_9(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_0 <= radians_load_node_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_1 <= wire_z_pipeff1_sub_result;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_1_w_q_range1421w(0) <= z_pipeff_1(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_10 <= z_pipenode_10_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_10_w_q_range8864w(0) <= z_pipeff_10(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_11 <= z_pipenode_11_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_11_w_q_range9666w(0) <= z_pipeff_11(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_12 <= z_pipenode_12_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_12_w_q_range10463w(0) <= z_pipeff_12(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_13 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_13 <= z_pipenode_13_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_2 <= z_pipenode_2_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_2_w_q_range2268w(0) <= z_pipeff_2(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_3 <= z_pipenode_3_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_3_w_q_range3110w(0) <= z_pipeff_3(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_4 <= z_pipenode_4_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_4_w_q_range3947w(0) <= z_pipeff_4(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_5 <= z_pipenode_5_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_5_w_q_range4779w(0) <= z_pipeff_5(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_6 <= z_pipenode_6_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_6_w_q_range5606w(0) <= z_pipeff_6(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_7 <= z_pipenode_7_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_7_w_q_range6428w(0) <= z_pipeff_7(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_8 <= z_pipenode_8_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_8_w_q_range7245w(0) <= z_pipeff_8(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_9 <= z_pipenode_9_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_9_w_q_range8057w(0) <= z_pipeff_9(33);
	wire_sincos_add_cin <= wire_sincosbitff_w_lg_w_q_range10746w10747w(0);
	sincos_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => wire_sincos_add_cin,
		dataa => delay_pipe_w,
		datab => post_estimate_w,
		result => wire_sincos_add_result
	  );
	x_pipenode_10_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_9(33),
		dataa => x_pipeff_9,
		datab => x_subnode_10_w,
		result => wire_x_pipenode_10_add_result
	  );
	x_pipenode_11_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_10(33),
		dataa => x_pipeff_10,
		datab => x_subnode_11_w,
		result => wire_x_pipenode_11_add_result
	  );
	x_pipenode_12_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_11(33),
		dataa => x_pipeff_11,
		datab => x_subnode_12_w,
		result => wire_x_pipenode_12_add_result
	  );
	x_pipenode_13_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_12(33),
		dataa => x_pipeff_12,
		datab => x_subnode_13_w,
		result => wire_x_pipenode_13_add_result
	  );
	x_pipenode_2_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_1(33),
		dataa => x_pipeff_1,
		datab => x_subnode_2_w,
		result => wire_x_pipenode_2_add_result
	  );
	x_pipenode_3_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_2(33),
		dataa => x_pipeff_2,
		datab => x_subnode_3_w,
		result => wire_x_pipenode_3_add_result
	  );
	x_pipenode_4_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_3(33),
		dataa => x_pipeff_3,
		datab => x_subnode_4_w,
		result => wire_x_pipenode_4_add_result
	  );
	x_pipenode_5_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_4(33),
		dataa => x_pipeff_4,
		datab => x_subnode_5_w,
		result => wire_x_pipenode_5_add_result
	  );
	x_pipenode_6_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_5(33),
		dataa => x_pipeff_5,
		datab => x_subnode_6_w,
		result => wire_x_pipenode_6_add_result
	  );
	x_pipenode_7_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_6(33),
		dataa => x_pipeff_6,
		datab => x_subnode_7_w,
		result => wire_x_pipenode_7_add_result
	  );
	x_pipenode_8_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_7(33),
		dataa => x_pipeff_7,
		datab => x_subnode_8_w,
		result => wire_x_pipenode_8_add_result
	  );
	x_pipenode_9_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_8(33),
		dataa => x_pipeff_8,
		datab => x_subnode_9_w,
		result => wire_x_pipenode_9_add_result
	  );
	y_pipeff1_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		dataa => y_pipeff_0,
		datab => y_subnode_1_w,
		result => wire_y_pipeff1_add_result
	  );
	y_pipenode_10_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_9(33),
		dataa => y_pipeff_9,
		datab => y_subnode_10_w,
		result => wire_y_pipenode_10_add_result
	  );
	y_pipenode_11_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_10(33),
		dataa => y_pipeff_10,
		datab => y_subnode_11_w,
		result => wire_y_pipenode_11_add_result
	  );
	y_pipenode_12_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_11(33),
		dataa => y_pipeff_11,
		datab => y_subnode_12_w,
		result => wire_y_pipenode_12_add_result
	  );
	y_pipenode_13_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_12(33),
		dataa => y_pipeff_12,
		datab => y_subnode_13_w,
		result => wire_y_pipenode_13_add_result
	  );
	y_pipenode_2_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_1(33),
		dataa => y_pipeff_1,
		datab => y_subnode_2_w,
		result => wire_y_pipenode_2_add_result
	  );
	y_pipenode_3_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_2(33),
		dataa => y_pipeff_2,
		datab => y_subnode_3_w,
		result => wire_y_pipenode_3_add_result
	  );
	y_pipenode_4_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_3(33),
		dataa => y_pipeff_3,
		datab => y_subnode_4_w,
		result => wire_y_pipenode_4_add_result
	  );
	y_pipenode_5_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_4(33),
		dataa => y_pipeff_4,
		datab => y_subnode_5_w,
		result => wire_y_pipenode_5_add_result
	  );
	y_pipenode_6_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_5(33),
		dataa => y_pipeff_5,
		datab => y_subnode_6_w,
		result => wire_y_pipenode_6_add_result
	  );
	y_pipenode_7_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_6(33),
		dataa => y_pipeff_6,
		datab => y_subnode_7_w,
		result => wire_y_pipenode_7_add_result
	  );
	y_pipenode_8_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_7(33),
		dataa => y_pipeff_7,
		datab => y_subnode_8_w,
		result => wire_y_pipenode_8_add_result
	  );
	y_pipenode_9_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_8(33),
		dataa => y_pipeff_8,
		datab => y_subnode_9_w,
		result => wire_y_pipenode_9_add_result
	  );
	z_pipeff1_sub :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		dataa => z_pipeff_0,
		datab => atannode_0_w,
		result => wire_z_pipeff1_sub_result
	  );
	z_pipenode_10_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_9(33),
		dataa => z_pipeff_9,
		datab => z_subnode_10_w,
		result => wire_z_pipenode_10_add_result
	  );
	z_pipenode_11_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_10(33),
		dataa => z_pipeff_10,
		datab => z_subnode_11_w,
		result => wire_z_pipenode_11_add_result
	  );
	z_pipenode_12_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_11(33),
		dataa => z_pipeff_11,
		datab => z_subnode_12_w,
		result => wire_z_pipenode_12_add_result
	  );
	z_pipenode_13_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_12(33),
		dataa => z_pipeff_12,
		datab => z_subnode_13_w,
		result => wire_z_pipenode_13_add_result
	  );
	z_pipenode_2_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_1(33),
		dataa => z_pipeff_1,
		datab => z_subnode_2_w,
		result => wire_z_pipenode_2_add_result
	  );
	z_pipenode_3_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_2(33),
		dataa => z_pipeff_2,
		datab => z_subnode_3_w,
		result => wire_z_pipenode_3_add_result
	  );
	z_pipenode_4_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_3(33),
		dataa => z_pipeff_3,
		datab => z_subnode_4_w,
		result => wire_z_pipenode_4_add_result
	  );
	z_pipenode_5_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_4(33),
		dataa => z_pipeff_4,
		datab => z_subnode_5_w,
		result => wire_z_pipenode_5_add_result
	  );
	z_pipenode_6_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_5(33),
		dataa => z_pipeff_5,
		datab => z_subnode_6_w,
		result => wire_z_pipenode_6_add_result
	  );
	z_pipenode_7_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_6(33),
		dataa => z_pipeff_6,
		datab => z_subnode_7_w,
		result => wire_z_pipenode_7_add_result
	  );
	z_pipenode_8_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_7(33),
		dataa => z_pipeff_7,
		datab => z_subnode_8_w,
		result => wire_z_pipenode_8_add_result
	  );
	z_pipenode_9_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_8(33),
		dataa => z_pipeff_8,
		datab => z_subnode_9_w,
		result => wire_z_pipenode_9_add_result
	  );
	cmx :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 3,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTHA => 34,
		LPM_WIDTHB => 34,
		LPM_WIDTHP => 68
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => multiplier_input_w,
		datab => z_pipeff_13,
		result => wire_cmx_result
	  );

 END RTL; --mysincos_altfp_sincos_cordic_m_a8e


--altfp_sincos_range CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" WIDTH_EXP=8 WIDTH_MAN=23 aclr circle clken clock data negcircle
--VERSION_BEGIN 13.0 cbx_altfp_sincos 2013:06:12:18:03:43:SJ cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_clshift 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END


--altfp_sincos_srrt CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" address basefraction incexponent incmantissa
--VERSION_BEGIN 13.0 cbx_altfp_sincos 2013:06:12:18:03:43:SJ cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_clshift 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.lpm_components.all;

--synthesis_resources = lpm_mux 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altfp_sincos_srrt_gra IS 
	 PORT 
	 ( 
		 address	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 basefraction	:	OUT  STD_LOGIC_VECTOR (35 DOWNTO 0);
		 incexponent	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 incmantissa	:	OUT  STD_LOGIC_VECTOR (55 DOWNTO 0)
	 ); 
 END mysincos_altfp_sincos_srrt_gra;

 ARCHITECTURE RTL OF mysincos_altfp_sincos_srrt_gra IS

	 SIGNAL  wire_mux2_data	:	STD_LOGIC_VECTOR (25599 DOWNTO 0);
	 SIGNAL  wire_mux2_data_2d	:	STD_LOGIC_2D(255 DOWNTO 0, 99 DOWNTO 0);
	 SIGNAL  wire_mux2_result	:	STD_LOGIC_VECTOR (99 DOWNTO 0);
 BEGIN

	basefraction <= wire_mux2_result(35 DOWNTO 0);
	incexponent <= wire_mux2_result(99 DOWNTO 92);
	incmantissa <= wire_mux2_result(91 DOWNTO 36);
	wire_mux2_data <= ( "00000000" & "10011010011011101110000001101101101100010100101011001000" & "00110110" & "1101100010100101011001100101" & "00000001" & "10011010011011101110000001101101101100010100101011010000" & "00011011" & "0110110001010010101100110010" & "00000000" & "10100110100110111011100000011011011011000101001010111000" & "00001101" & "1011011000101001010110011001" & "00000001" & "10100110100110111011100000011011011011000101001010110000" & "00000110" & "1101101100010100101011001101" & "00000000" & "10101001101001101110111000000110110110110001010010110000" & "00000011" & "0110110110001010010101100110" & "00000000" & "11010100110100110111011100000011011011011000101001100000" & "10000001" & "1011011011000101001010110011" & "00000000" & "11101010011010011011101110000001101101101100010100011000" & "11000000" & "1101101101100010100101011010" & "00000000" & "11110101001101001101110111000000110110110110001010011000" & "11100000" & "0110110110110001010010101101" & "00000000" & "11111010100110100110111011100000011011011011000101010000" & "01110000" & "0011011011011000101001010110" & "00000001" & "11111010100110100110111011100000011011011011000101010000" & "10111000" & "0001101101101100010100101011" & "00000010" & "11111010100110100110111011100000011011011011000101010000" & "11011100" & "0000110110110110001010010110" & "00000011" & "11111010100110100110111011100000011011011011000100101000" & "11101110" & "0000011011011011000101001011" & "00000000" & "10001111101010011010011011101110000001101101101100011000" & "01110111" & "0000001101101101100010100101" & "00000001" & "10001111101010011010011011101110000001101101101100100000" & "10111011" & "1000000110110110110001010011" & "00000000" & "10100011111010100110100110111011100000011011011011001000" & "11011101" & "1100000011011011011000101001" & "00000000" & "11010001111101010011010011011101110000001101101101010000" & "01101110" & "1110000001101101101100010101" & "00000000" & "11101000111110101001101001101110111000000110110110111000" & "00110111" & "0111000000110110110110001010"
 & "00000000" & "11110100011111010100110100110111011100000011011011011000" & "10011011" & "1011100000011011011011000101" & "00000000" & "11111010001111101010011010011011101110000001101101101000" & "01001101" & "1101110000001101101101100011" & "00000001" & "11111010001111101010011010011011101110000001101110000000" & "10100110" & "1110111000000110110110110001" & "00000000" & "10111110100011111010100110100110111011100000011011100000" & "11010011" & "0111011100000011011011011001" & "00000001" & "10111110100011111010100110100110111011100000011011101000" & "01101001" & "1011101110000001101101101100" & "00000000" & "10101111101000111110101001101001101110111000000110111000" & "00110100" & "1101110111000000110110110110" & "00000001" & "10101111101000111110101001101001101110111000000110110000" & "10011010" & "0110111011100000011011011011" & "00000000" & "10101011111010001111101010011010011011101110000001110000" & "01001101" & "0011011101110000001101101110" & "00000000" & "11010101111101000111110101001101001101110111000000111000" & "10100110" & "1001101110111000000110110111" & "00000000" & "11101010111110100011111010100110100110111011100000110000" & "01010011" & "0100110111011100000011011011" & "00000001" & "11101010111110100011111010100110100110111011100000100000" & "10101001" & "1010011011101110000001101110" & "00000010" & "11101010111110100011111010100110100110111011011111111000" & "11010100" & "1101001101110111000000110111" & "00000000" & "10011101010111110100011111010100110100110111011100000000" & "11101010" & "0110100110111011100000011011" & "00000001" & "10011101010111110100011111010100110100110111011100011000" & "11110101" & "0011010011011101110000001110" & "00000010" & "10011101010111110100011111010100110100110111011100011000" & "11111010" & "1001101001101110111000000111" & "00000011" & "10011101010111110100011111010100110100110111011100011000" & "01111101" & "0100110100110111011100000011" & "00000100" & "10011101010111110100011111010100110100110111011110010000" & "00111110" & "1010011010011011101110000010" & "00000000"
 & "10000100111010101111101000111110101001101001101111000000" & "00011111" & "0101001101001101110111000001" & "00000000" & "11000010011101010111110100011111010100110100110111011000" & "10001111" & "1010100110100110111011100000" & "00000000" & "11100001001110101011111010001111101010011010011011110000" & "01000111" & "1101010011010011011101110000" & "00000000" & "11110000100111010101111101000111110101001101001110000000" & "10100011" & "1110101001101001101110111000" & "00000000" & "11111000010011101010111110100011111010100110100110111000" & "11010001" & "1111010100110100110111011100" & "00000000" & "11111100001001110101011111010001111101010011010011011000" & "11101000" & "1111101010011010011011101110" & "00000000" & "11111110000100111010101111101000111110101001101001110000" & "11110100" & "0111110101001101001101110111" & "00000001" & "11111110000100111010101111101000111110101001101010000000" & "11111010" & "0011111010100110100110111100" & "00000010" & "11111110000100111010101111101000111110101001101001110000" & "01111101" & "0001111101010011010011011110" & "00000000" & "10011111110000100111010101111101000111110101001101011000" & "10111110" & "1000111110101001101001101111" & "00000001" & "10011111110000100111010101111101000111110101001101100000" & "01011111" & "0100011111010100110100110111" & "00000000" & "10100111111100001001110101011111010001111101010011010000" & "10101111" & "1010001111101010011010011100" & "00000001" & "10100111111100001001110101011111010001111101010011100000" & "01010111" & "1101000111110101001101001110" & "00000010" & "10100111111100001001110101011111010001111101010011010000" & "10101011" & "1110100011111010100110100111" & "00000000" & "10010100111111100001001110101011111010001111101010011000" & "11010101" & "1111010001111101010011010011" & "00000001" & "10010100111111100001001110101011111010001111101010101000" & "11101010" & "1111101000111110101001101010" & "00000000" & "10100101001111111000010011101010111110100011111010101000" & "01110101" & "0111110100011111010100110101" & "00000001" & "10100101001111111000010011101010111110100011111010101000"
 & "00111010" & "1011111010001111101010011010" & "00000000" & "10101001010011111110000100111010101111101000111110101000" & "10011101" & "0101111101000111110101001101" & "00000001" & "10101001010011111110000100111010101111101000111110111000" & "01001110" & "1010111110100011111010100111" & "00000010" & "10101001010011111110000100111010101111101000111110111000" & "00100111" & "0101011111010001111101010011" & "00000011" & "10101001010011111110000100111010101111101000111110111000" & "00010011" & "1010101111101000111110101010" & "00000100" & "10101001010011111110000100111010101111101000111110111000" & "00001001" & "1101010111110100011111010101" & "00000101" & "10101001010011111110000100111010101111101001000000110000" & "10000100" & "1110101011111010001111101010" & "00000000" & "10000010101001010011111110000100111010101111101001001000" & "11000010" & "0111010101111101000111110101" & "00000001" & "10000010101001010011111110000100111010101111101001010000" & "11100001" & "0011101010111110100011111011" & "00000010" & "10000010101001010011111110000100111010101111101000111000" & "11110000" & "1001110101011111010001111101" & "00000011" & "10000010101001010011111110000100111010101111101001100000" & "11111000" & "0100111010101111101000111111" & "00000000" & "10001000001010100101001111111000010011101010111110100000" & "11111100" & "0010011101010111110100011111" & "00000001" & "10001000001010100101001111111000010011101010111110100000" & "11111110" & "0001001110101011111010010000" & "00000010" & "10001000001010100101001111111000010011101010111110100000" & "01111111" & "0000100111010101111101001000" & "00000000" & "10010001000001010100101001111111000010011101011000010000" & "00111111" & "1000010011101010111110100100" & "00000000" & "11001000100000101010010100111111100001001110101011111000" & "10011111" & "1100001001110101011111010010" & "00000000" & "11100100010000010101001010011111110000100111010101111000" & "01001111" & "1110000100111010101111101001" & "00000001" & "11100100010000010101001010011111110000100111010101110000" & "10100111"
 & "1111000010011101010111110100" & "00000010" & "11100100010000010101001010011111110000100111010110001000" & "01010011" & "1111100001001110101011111010" & "00000000" & "10011100100010000010101001010011111110000100111010111000" & "00101001" & "1111110000100111010101111101" & "00000001" & "10011100100010000010101001010011111110000100111010111000" & "10010100" & "1111111000010011101010111111" & "00000010" & "10011100100010000010101001010011111110000100111010110000" & "01001010" & "0111111100001001110101011111" & "00000000" & "10010011100100010000010101001010011111110000100111011000" & "10100101" & "0011111110000100111010110000" & "00000000" & "11001001110010001000001010100101001111111000010011101000" & "01010010" & "1001111111000010011101011000" & "00000000" & "11100100111001000100000101010010100111111100001001111000" & "10101001" & "0100111111100001001110101100" & "00000001" & "11100100111001000100000101010010100111111100001001101000" & "01010100" & "1010011111110000100111010110" & "00000000" & "10111001001110010001000001010100101001111111000010011000" & "00101010" & "0101001111111000010011101011" & "00000000" & "11011100100111001000100000101010010100111111100001011000" & "00010101" & "0010100111111100001001110101" & "00000001" & "11011100100111001000100000101010010100111111100001011000" & "00001010" & "1001010011111110000100111011" & "00000000" & "10110111001001110010001000001010100101001111111000011000" & "00000101" & "0100101001111111000010011101" & "00000000" & "11011011100100111001000100000101010010100111111100001000" & "10000010" & "1010010100111111100001001111" & "00000001" & "11011011100100111001000100000101010010100111111011111000" & "01000001" & "0101001010011111110000100111" & "00000010" & "11011011100100111001000100000101010010100111111100001000" & "00100000" & "1010100101001111111000010100" & "00000011" & "11011011100100111001000100000101010010100111111100100000" & "00010000" & "0101010010100111111100001010" & "00000100" & "11011011100100111001000100000101010010100111111010111000" & "10001000" & "0010101001010011111110000101"
 & "00000101" & "11011011100100111001000100000101010010100111111001101000" & "01000100" & "0001010100101001111111000010" & "00000000" & "10000011011011100100111001000100000101010010101000000000" & "00100010" & "0000101010010100111111100001" & "00000000" & "11000001101101110010011100100010000010101001010100001000" & "10010001" & "0000010101001010011111110001" & "00000001" & "11000001101101110010011100100010000010101001010011110000" & "11001000" & "1000001010100101001111111000" & "00000010" & "11000001101101110010011100100010000010101001010100001000" & "11100100" & "0100000101010010100111111100" & "00000000" & "10011000001101101110010011100100010000010101001010100000" & "01110010" & "0010000010101001010011111110" & "00000000" & "11001100000110110111001001110010001000001010100101010000" & "00111001" & "0001000001010100101001111111" & "00000000" & "11100110000011011011100100111001000100000101010010101000" & "10011100" & "1000100000101010010101000000" & "00000000" & "11110011000001101101110010011100100010000010101001001000" & "01001110" & "0100010000010101001010100000" & "00000000" & "11111001100000110110111001001110010001000001010100101000" & "00100111" & "0010001000001010100101010000" & "00000001" & "11111001100000110110111001001110010001000001010100101000" & "10010011" & "1001000100000101010010101000" & "00000000" & "10111110011000001101101110010011100100010000010101010000" & "11001001" & "1100100010000010101001010100" & "00000001" & "10111110011000001101101110010011100100010000010101011000" & "11100100" & "1110010001000001010100101010" & "00000010" & "10111110011000001101101110010011100100010000010101000000" & "01110010" & "0111001000100000101010010101" & "00000011" & "10111110011000001101101110010011100100010000010101110000" & "10111001" & "0011100100010000010101001010" & "00000000" & "10001011111001100000110110111001001110010001000001011000" & "11011100" & "1001110010001000001010100101" & "00000001" & "10001011111001100000110110111001001110010001000001010000" & "01101110" & "0100111001000100000101010011" & "00000000"
 & "10100010111110011000001101101110010011100100010000010000" & "10110111" & "0010011100100010000010101001" & "00000001" & "10100010111110011000001101101110010011100100010000011000" & "11011011" & "1001001110010001000001010101" & "00000010" & "10100010111110011000001101101110010011100100010000011000" & "01101101" & "1100100111001000100000101010" & "00000011" & "10100010111110011000001101101110010011100100010000011000" & "00110110" & "1110010011100100010000010101" & "00000100" & "10100010111110011000001101101110010011100100010000011000" & "00011011" & "0111001001110010001000001011" & "00000101" & "10100010111110011000001101101110010011100100010000011000" & "00001101" & "1011100100111001000100000101" & "00000110" & "10100010111110011000001101101110010011100100010000011000" & "00000110" & "1101110010011100100010000011" & "00000111" & "10100010111110011000001101101110010011100100010000011000" & "10000011" & "0110111001001110010001000001" & "00001000" & "10100010111110011000001101101110010011100101100001111000" & "11000001" & "1011011100100111001000100001" & "00001001" & "10100010111110011000001101101110010011100100010000011000" & "01100000" & "1101101110010011100100010000" & "00001010" & "10100010111110011000001101101110010011100100010000011000" & "00110000" & "0110110111001001110010001000" & "00001011" & "10100010111110011000001101101110010011100100010000011000" & "10011000" & "0011011011100100111001000100" & "00001100" & "10100010111110011000001101101110010011100100010000011000" & "11001100" & "0001101101110010011100100010" & "00001101" & "10100010111110011000001101101110010011100100010000011000" & "11100110" & "0000110110111001001110010001" & "00001110" & "10100010111110011000001101101110010011100100010000011000" & "11110011" & "0000011011011100100111001001" & "00001111" & "10100010111110011000001101101110010011100100010000011000" & "11111001" & "1000001101101110010011100100" & "00010000" & "10100010111110011000001101101110010011100100010000011000" & "01111100" & "1100000110110111001001110010" & "00010001" & "10100010111110011000001101101110001001011000010110111000"
 & "10111110" & "0110000011011011100100111001" & "00010010" & "10100010111110011000001101101110010011100100010000011000" & "01011111" & "0011000001101101110010011101" & "00010011" & "10100010111110011000001101101110011000101010001101001000" & "00101111" & "1001100000110110111001001110" & "00010100" & "10100010111110011000001101101110010011100100010000011000" & "00010111" & "1100110000011011011100100111" & "00010101" & "10100010111110011000001101101110010011100100010000011000" & "10001011" & "1110011000001101101110010100" & "00010110" & "10100010111110011000001101101110010011100100010000011000" & "01000101" & "1111001100000110110111001010" & "00010111" & "10100010111110011000001101101110010011100100010000011000" & "10100010" & "1111100110000011011011100101" & "00011000" & "10100010111110011000001101110000110110100010101000101000" & "01010001" & "0111110011000001101101110010" & "00011001" & "10100010111110011000001101101110010011100100010000011000" & "00101000" & "1011111001100000110110111001" & "00011010" & "10100010111110011000001101101110010011100100010000011000" & "00010100" & "0101111100110000011011011101" & "00011011" & "10100010111110011000001101101110010011100100010000011000" & "00001010" & "0010111110011000001101101110" & "00011100" & "10100010111110011000001101101110010011100100010000011000" & "00000101" & "0001011111001100000110110111" & "00011101" & "10100010111110011000001101101110010011100100010000011000" & "00000010" & "1000101111100110000011011100" & "00011110" & "10100010111110011000001101101110010011100100010000011000" & "00000001" & "0100010111110011000001101110" & "00011111" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "1010001011111001100000110111" & "00100000" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0101000101111100110000011011" & "00100001" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0010100010111110011000001110" & "00100010" & "10100010111110011000001101101110010011100100010000011000" & "00000000"
 & "0001010001011111001100000111" & "00100011" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000101000101111100110000011" & "00100100" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000010100010111110011000010" & "00100101" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000001010001011111001100001" & "00100110" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000000101000101111100110000" & "00100111" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000000010100010111110011000" & "00101000" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000000001010001011111001100" & "00101001" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000000000101000101111100110" & "00101010" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000000000010100010111110011" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
	loop36 : FOR i IN 0 TO 255 GENERATE
		loop37 : FOR j IN 0 TO 99 GENERATE
			wire_mux2_data_2d(i, j) <= wire_mux2_data(i*100+j);
		END GENERATE loop37;
	END GENERATE loop36;
	mux2 :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 256,
		LPM_WIDTH => 100,
		LPM_WIDTHS => 8
	  )
	  PORT MAP ( 
		data => wire_mux2_data_2d,
		result => wire_mux2_result,
		sel => address
	  );

 END RTL; --mysincos_altfp_sincos_srrt_gra


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" WIDTH=32 WIDTHAD=5 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=16 WIDTHAD=4 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altpriority_encoder_3e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END mysincos_altpriority_encoder_3e8;

 ARCHITECTURE RTL OF mysincos_altpriority_encoder_3e8 IS

 BEGIN

	q(0) <= ( data(1));
	zero <= (NOT (data(0) OR data(1)));

 END RTL; --mysincos_altpriority_encoder_3e8


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altpriority_encoder_3v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0)
	 ); 
 END mysincos_altpriority_encoder_3v7;

 ARCHITECTURE RTL OF mysincos_altpriority_encoder_3v7 IS

 BEGIN

	q(0) <= ( data(1));

 END RTL; --mysincos_altpriority_encoder_3v7

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altpriority_encoder_6v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0)
	 ); 
 END mysincos_altpriority_encoder_6v7;

 ARCHITECTURE RTL OF mysincos_altpriority_encoder_6v7 IS

	 SIGNAL  wire_altpriority_encoder10_w_lg_w_lg_zero13017w13018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_zero13019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_zero13017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_w_lg_zero13019w13020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder9_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  mysincos_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  mysincos_altpriority_encoder_3v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder10_w_lg_zero13017w & wire_altpriority_encoder10_w_lg_w_lg_zero13019w13020w);
	wire_altpriority_encoder10_w_lg_w_lg_zero13017w13018w(0) <= wire_altpriority_encoder10_w_lg_zero13017w(0) AND wire_altpriority_encoder10_q(0);
	wire_altpriority_encoder10_w_lg_zero13019w(0) <= wire_altpriority_encoder10_zero AND wire_altpriority_encoder9_q(0);
	wire_altpriority_encoder10_w_lg_zero13017w(0) <= NOT wire_altpriority_encoder10_zero;
	wire_altpriority_encoder10_w_lg_w_lg_zero13019w13020w(0) <= wire_altpriority_encoder10_w_lg_zero13019w(0) OR wire_altpriority_encoder10_w_lg_w_lg_zero13017w13018w(0);
	altpriority_encoder10 :  mysincos_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder10_q,
		zero => wire_altpriority_encoder10_zero
	  );
	altpriority_encoder9 :  mysincos_altpriority_encoder_3v7
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder9_q
	  );

 END RTL; --mysincos_altpriority_encoder_6v7


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altpriority_encoder_6e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END mysincos_altpriority_encoder_6e8;

 ARCHITECTURE RTL OF mysincos_altpriority_encoder_6e8 IS

	 SIGNAL  wire_altpriority_encoder11_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder12_w_lg_w_lg_zero13035w13036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_zero13037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_zero13035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_w_lg_zero13037w13038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_zero	:	STD_LOGIC;
	 COMPONENT  mysincos_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder12_w_lg_zero13035w & wire_altpriority_encoder12_w_lg_w_lg_zero13037w13038w);
	zero <= (wire_altpriority_encoder11_zero AND wire_altpriority_encoder12_zero);
	altpriority_encoder11 :  mysincos_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder11_q,
		zero => wire_altpriority_encoder11_zero
	  );
	wire_altpriority_encoder12_w_lg_w_lg_zero13035w13036w(0) <= wire_altpriority_encoder12_w_lg_zero13035w(0) AND wire_altpriority_encoder12_q(0);
	wire_altpriority_encoder12_w_lg_zero13037w(0) <= wire_altpriority_encoder12_zero AND wire_altpriority_encoder11_q(0);
	wire_altpriority_encoder12_w_lg_zero13035w(0) <= NOT wire_altpriority_encoder12_zero;
	wire_altpriority_encoder12_w_lg_w_lg_zero13037w13038w(0) <= wire_altpriority_encoder12_w_lg_zero13037w(0) OR wire_altpriority_encoder12_w_lg_w_lg_zero13035w13036w(0);
	altpriority_encoder12 :  mysincos_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder12_q,
		zero => wire_altpriority_encoder12_zero
	  );

 END RTL; --mysincos_altpriority_encoder_6e8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altpriority_encoder_bv7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0)
	 ); 
 END mysincos_altpriority_encoder_bv7;

 ARCHITECTURE RTL OF mysincos_altpriority_encoder_bv7 IS

	 SIGNAL  wire_altpriority_encoder7_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_w_lg_w_lg_zero13008w13009w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_w_lg_zero13010w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_w_lg_zero13008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_w_lg_w_lg_zero13010w13011w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_zero	:	STD_LOGIC;
	 COMPONENT  mysincos_altpriority_encoder_6v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  mysincos_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder8_w_lg_zero13008w & wire_altpriority_encoder8_w_lg_w_lg_zero13010w13011w);
	altpriority_encoder7 :  mysincos_altpriority_encoder_6v7
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder7_q
	  );
	loop38 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder8_w_lg_w_lg_zero13008w13009w(i) <= wire_altpriority_encoder8_w_lg_zero13008w(0) AND wire_altpriority_encoder8_q(i);
	END GENERATE loop38;
	loop39 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder8_w_lg_zero13010w(i) <= wire_altpriority_encoder8_zero AND wire_altpriority_encoder7_q(i);
	END GENERATE loop39;
	wire_altpriority_encoder8_w_lg_zero13008w(0) <= NOT wire_altpriority_encoder8_zero;
	loop40 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder8_w_lg_w_lg_zero13010w13011w(i) <= wire_altpriority_encoder8_w_lg_zero13010w(i) OR wire_altpriority_encoder8_w_lg_w_lg_zero13008w13009w(i);
	END GENERATE loop40;
	altpriority_encoder8 :  mysincos_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder8_q,
		zero => wire_altpriority_encoder8_zero
	  );

 END RTL; --mysincos_altpriority_encoder_bv7


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altpriority_encoder_be8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END mysincos_altpriority_encoder_be8;

 ARCHITECTURE RTL OF mysincos_altpriority_encoder_be8 IS

	 SIGNAL  wire_altpriority_encoder13_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder14_w_lg_w_lg_zero13045w13046w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_zero13047w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_zero13045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_w_lg_zero13047w13048w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_zero	:	STD_LOGIC;
	 COMPONENT  mysincos_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder14_w_lg_zero13045w & wire_altpriority_encoder14_w_lg_w_lg_zero13047w13048w);
	zero <= (wire_altpriority_encoder13_zero AND wire_altpriority_encoder14_zero);
	altpriority_encoder13 :  mysincos_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder13_q,
		zero => wire_altpriority_encoder13_zero
	  );
	loop41 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder14_w_lg_w_lg_zero13045w13046w(i) <= wire_altpriority_encoder14_w_lg_zero13045w(0) AND wire_altpriority_encoder14_q(i);
	END GENERATE loop41;
	loop42 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder14_w_lg_zero13047w(i) <= wire_altpriority_encoder14_zero AND wire_altpriority_encoder13_q(i);
	END GENERATE loop42;
	wire_altpriority_encoder14_w_lg_zero13045w(0) <= NOT wire_altpriority_encoder14_zero;
	loop43 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder14_w_lg_w_lg_zero13047w13048w(i) <= wire_altpriority_encoder14_w_lg_zero13047w(i) OR wire_altpriority_encoder14_w_lg_w_lg_zero13045w13046w(i);
	END GENERATE loop43;
	altpriority_encoder14 :  mysincos_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder14_q,
		zero => wire_altpriority_encoder14_zero
	  );

 END RTL; --mysincos_altpriority_encoder_be8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altpriority_encoder_r08 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0)
	 ); 
 END mysincos_altpriority_encoder_r08;

 ARCHITECTURE RTL OF mysincos_altpriority_encoder_r08 IS

	 SIGNAL  wire_altpriority_encoder5_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder6_w_lg_w_lg_zero12999w13000w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder6_w_lg_zero13001w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder6_w_lg_zero12999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder6_w_lg_w_lg_zero13001w13002w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder6_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder6_zero	:	STD_LOGIC;
	 COMPONENT  mysincos_altpriority_encoder_bv7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  mysincos_altpriority_encoder_be8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder6_w_lg_zero12999w & wire_altpriority_encoder6_w_lg_w_lg_zero13001w13002w);
	altpriority_encoder5 :  mysincos_altpriority_encoder_bv7
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder5_q
	  );
	loop44 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder6_w_lg_w_lg_zero12999w13000w(i) <= wire_altpriority_encoder6_w_lg_zero12999w(0) AND wire_altpriority_encoder6_q(i);
	END GENERATE loop44;
	loop45 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder6_w_lg_zero13001w(i) <= wire_altpriority_encoder6_zero AND wire_altpriority_encoder5_q(i);
	END GENERATE loop45;
	wire_altpriority_encoder6_w_lg_zero12999w(0) <= NOT wire_altpriority_encoder6_zero;
	loop46 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder6_w_lg_w_lg_zero13001w13002w(i) <= wire_altpriority_encoder6_w_lg_zero13001w(i) OR wire_altpriority_encoder6_w_lg_w_lg_zero12999w13000w(i);
	END GENERATE loop46;
	altpriority_encoder6 :  mysincos_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder6_q,
		zero => wire_altpriority_encoder6_zero
	  );

 END RTL; --mysincos_altpriority_encoder_r08


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=16 WIDTHAD=4 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altpriority_encoder_rf8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END mysincos_altpriority_encoder_rf8;

 ARCHITECTURE RTL OF mysincos_altpriority_encoder_rf8 IS

	 SIGNAL  wire_altpriority_encoder15_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder16_w_lg_w_lg_zero13055w13056w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_zero13057w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_zero13055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_w_lg_zero13057w13058w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_zero	:	STD_LOGIC;
	 COMPONENT  mysincos_altpriority_encoder_be8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder16_w_lg_zero13055w & wire_altpriority_encoder16_w_lg_w_lg_zero13057w13058w);
	zero <= (wire_altpriority_encoder15_zero AND wire_altpriority_encoder16_zero);
	altpriority_encoder15 :  mysincos_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder15_q,
		zero => wire_altpriority_encoder15_zero
	  );
	loop47 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder16_w_lg_w_lg_zero13055w13056w(i) <= wire_altpriority_encoder16_w_lg_zero13055w(0) AND wire_altpriority_encoder16_q(i);
	END GENERATE loop47;
	loop48 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder16_w_lg_zero13057w(i) <= wire_altpriority_encoder16_zero AND wire_altpriority_encoder15_q(i);
	END GENERATE loop48;
	wire_altpriority_encoder16_w_lg_zero13055w(0) <= NOT wire_altpriority_encoder16_zero;
	loop49 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder16_w_lg_w_lg_zero13057w13058w(i) <= wire_altpriority_encoder16_w_lg_zero13057w(i) OR wire_altpriority_encoder16_w_lg_w_lg_zero13055w13056w(i);
	END GENERATE loop49;
	altpriority_encoder16 :  mysincos_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder16_q,
		zero => wire_altpriority_encoder16_zero
	  );

 END RTL; --mysincos_altpriority_encoder_rf8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altpriority_encoder_qb6 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0)
	 ); 
 END mysincos_altpriority_encoder_qb6;

 ARCHITECTURE RTL OF mysincos_altpriority_encoder_qb6 IS

	 SIGNAL  wire_altpriority_encoder3_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder4_w_lg_w_lg_zero12990w12991w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder4_w_lg_zero12992w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder4_w_lg_zero12990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder4_w_lg_w_lg_zero12992w12993w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder4_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder4_zero	:	STD_LOGIC;
	 COMPONENT  mysincos_altpriority_encoder_r08
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  mysincos_altpriority_encoder_rf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder4_w_lg_zero12990w & wire_altpriority_encoder4_w_lg_w_lg_zero12992w12993w);
	altpriority_encoder3 :  mysincos_altpriority_encoder_r08
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder3_q
	  );
	loop50 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder4_w_lg_w_lg_zero12990w12991w(i) <= wire_altpriority_encoder4_w_lg_zero12990w(0) AND wire_altpriority_encoder4_q(i);
	END GENERATE loop50;
	loop51 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder4_w_lg_zero12992w(i) <= wire_altpriority_encoder4_zero AND wire_altpriority_encoder3_q(i);
	END GENERATE loop51;
	wire_altpriority_encoder4_w_lg_zero12990w(0) <= NOT wire_altpriority_encoder4_zero;
	loop52 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder4_w_lg_w_lg_zero12992w12993w(i) <= wire_altpriority_encoder4_w_lg_zero12992w(i) OR wire_altpriority_encoder4_w_lg_w_lg_zero12990w12991w(i);
	END GENERATE loop52;
	altpriority_encoder4 :  mysincos_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder4_q,
		zero => wire_altpriority_encoder4_zero
	  );

 END RTL; --mysincos_altpriority_encoder_qb6

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 8 lpm_clshift 2 lpm_mult 1 lpm_mux 1 reg 780 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altfp_sincos_range_79c IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 circle	:	OUT  STD_LOGIC_VECTOR (35 DOWNTO 0);
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
		 negcircle	:	OUT  STD_LOGIC_VECTOR (35 DOWNTO 0)
	 ); 
 END mysincos_altfp_sincos_range_79c;

 ARCHITECTURE RTL OF mysincos_altfp_sincos_range_79c IS

	 SIGNAL  wire_fp_range_table1_basefraction	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_fp_range_table1_incexponent	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_fp_range_table1_incmantissa	:	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  wire_clz23_data	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_clz23_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL	 basefractiondelff	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 basefractionff	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cbfd_0	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cbfd_1	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cbfd_2	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cbfd_3	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cbfd_4	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cbfd_5	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 circleff	:	STD_LOGIC_VECTOR(36 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exponentff	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 incexponentff	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 incmantissaff	:	STD_LOGIC_VECTOR(55 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 leadff	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mantissadelff	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mantissaff	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mantissamultiplierff	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 multipliernormff	:	STD_LOGIC_VECTOR(77 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 negbasefractiondelff	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 negcircleff	:	STD_LOGIC_VECTOR(36 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 negrangeexponentff4	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 negrangeexponentff5	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_negrangeexponentff5_w_lg_w_lg_w_q_range11460w11464w11465w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_negrangeexponentff5_w_lg_w_q_range11460w11462w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_negrangeexponentff5_w_lg_w_q_range11460w11464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_negrangeexponentff5_w_q_range11461w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_negrangeexponentff5_w_q_range11460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rangeexponentff_0	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rangeexponentff_1	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rangeexponentff_2	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rangeexponentff_3	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rangeexponentff_4	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rangeexponentff_5	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rangeexponentff_5_w_q_range11463w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL	 rotateff	:	STD_LOGIC_VECTOR(77 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rotateff_w_lg_w_q_range11477w11479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11481w11483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11484w11486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11487w11489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11490w11492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11493w11495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11496w11498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11499w11501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11502w11504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11505w11507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11508w11510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11511w11513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11514w11516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11517w11519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11520w11522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11523w11525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11526w11528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11529w11531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11532w11534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11535w11537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11538w11540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11541w11543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11544w11546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11547w11549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11550w11552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11553w11555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11556w11558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11559w11561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11562w11564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11565w11567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11568w11570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11571w11573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11574w11576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11577w11579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11580w11582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11583w11585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 tableaddressff	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_circle_add_dataa	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_circle_add_datab	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_circle_add_result	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_exponent_adjust_sub_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_exponent_adjust_sub_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_negbasedractiondel_sub_dataa	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_negbasedractiondel_sub_result	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_negcircle_add_dataa	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_negcircle_add_datab	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_negcircle_add_result	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_negrangeexponent_sub4_dataa	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_negrangeexponent_sub4_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_negrangeexponent_sub5_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_negrangeexponent_sub5_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_rangeexponent_sub1_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_rangeexponent_sub1_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_rangeexponent_sub5_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_rangeexponent_sub5_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_csftin_result	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_fp_lsft_rsft78_distance	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_negrangeexponentff5_w_lg_w_lg_w_lg_w_q_range11460w11464w11465w11466w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_fp_lsft_rsft78_result	:	STD_LOGIC_VECTOR (77 DOWNTO 0);
	 SIGNAL  wire_mult23x56_result	:	STD_LOGIC_VECTOR (78 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11069w11072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11116w11123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11116w11119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11121w11128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11121w11124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11126w11133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11126w11129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11131w11138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11131w11134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11136w11143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11136w11139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11141w11148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11141w11144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11146w11153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11146w11149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11151w11158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11151w11154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11156w11163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11156w11159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11161w11168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11161w11164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11070w11078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11070w11073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11166w11173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11166w11169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11171w11178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11171w11174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11176w11183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11176w11179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11181w11188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11181w11184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11186w11193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11186w11189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11191w11198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11191w11194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11196w11203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11196w11199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11201w11208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11201w11204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11206w11213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11206w11209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11211w11218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11211w11214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11076w11083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11076w11079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11216w11223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11216w11219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11221w11228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11221w11224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11226w11233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11226w11229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11231w11238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11231w11234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11236w11243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11236w11239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11241w11248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11241w11244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11246w11253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11246w11249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11251w11258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11251w11254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11256w11263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11256w11259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11261w11268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11261w11264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11081w11088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11081w11084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11266w11273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11266w11269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11271w11278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11271w11274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11276w11283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11276w11279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11281w11288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11281w11284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11286w11293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11286w11289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11291w11298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11291w11294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11296w11303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11296w11299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11301w11308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11301w11304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11306w11313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11306w11309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11311w11318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11311w11314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11086w11093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11086w11089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11316w11323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11316w11319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11321w11328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11321w11324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11326w11333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11326w11329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11331w11338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11331w11334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11336w11343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11336w11339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11341w11348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11341w11344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11346w11353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11346w11349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11351w11358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11351w11354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11356w11363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11356w11359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11361w11368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11361w11364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11091w11098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11091w11094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11366w11373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11366w11369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11371w11378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11371w11374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11376w11383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11376w11379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11381w11388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11381w11384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11386w11393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11386w11389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11391w11398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11391w11394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11396w11403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11396w11399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11401w11408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11401w11404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11406w11413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11406w11409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11411w11418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11411w11414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11096w11103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11096w11099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11416w11423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11416w11419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11421w11428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11421w11424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11426w11433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11426w11429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11431w11438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11431w11434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11436w11443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11436w11439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11441w11448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11441w11444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11446w11453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11446w11449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11451w11457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11451w11454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11101w11108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11101w11104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11106w11113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11106w11109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11111w11118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11111w11114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  basefractiondelnode_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  basefractionnode_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  circlenode_w :	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  const_23_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  incexponentnode_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  incmantissanode_w :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  leadnode_w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  mantissaexponentnode_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  mantissamultipliernode_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  multipliernode_w :	STD_LOGIC_VECTOR (78 DOWNTO 0);
	 SIGNAL  multipliernormnode_w :	STD_LOGIC_VECTOR (77 DOWNTO 0);
	 SIGNAL  negbasefractiondelnode_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  negcirclenode_w :	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  negrotatenode_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  rotatenode_w :	STD_LOGIC_VECTOR (77 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_data_range11039w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_data_range11040w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  mysincos_altfp_sincos_srrt_gra
	 PORT
	 ( 
		address	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		basefraction	:	OUT  STD_LOGIC_VECTOR(35 DOWNTO 0);
		incexponent	:	OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		incmantissa	:	OUT  STD_LOGIC_VECTOR(55 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  mysincos_altpriority_encoder_qb6
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_clshift
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_SHIFTTYPE	:	STRING := "LOGICAL";
		LPM_WIDTH	:	NATURAL;
		LPM_WIDTHDIST	:	NATURAL;
		lpm_type	:	STRING := "lpm_clshift"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		direction	:	IN STD_LOGIC := '0';
		distance	:	IN STD_LOGIC_VECTOR(LPM_WIDTHDIST-1 DOWNTO 0);
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		underflow	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_mult
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTHA	:	NATURAL;
		LPM_WIDTHB	:	NATURAL;
		LPM_WIDTHP	:	NATURAL;
		LPM_WIDTHS	:	NATURAL := 1;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_mult"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTHA-1 DOWNTO 0);
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTHB-1 DOWNTO 0);
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHP-1 DOWNTO 0);
		sum	:	IN STD_LOGIC_VECTOR(LPM_WIDTHS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11069w11072w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11069w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11116w11123w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11116w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11116w11119w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11116w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11121w11128w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11121w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11121w11124w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11121w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11126w11133w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11126w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11126w11129w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11126w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11131w11138w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11131w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11131w11134w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11131w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11136w11143w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11136w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11136w11139w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11136w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11141w11148w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11141w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11141w11144w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11141w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11146w11153w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11146w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11146w11149w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11146w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11151w11158w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11151w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11151w11154w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11151w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11156w11163w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11156w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11156w11159w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11156w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11161w11168w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11161w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11161w11164w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11161w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11070w11078w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11070w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11070w11073w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11070w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11166w11173w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11166w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11166w11169w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11166w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11171w11178w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11171w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11171w11174w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11171w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11176w11183w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11176w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11176w11179w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11176w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11181w11188w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11181w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11181w11184w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11181w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11186w11193w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11186w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11186w11189w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11186w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11191w11198w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11191w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11191w11194w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11191w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11196w11203w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11196w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11196w11199w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11196w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11201w11208w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11201w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11201w11204w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11201w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11206w11213w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11206w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11206w11209w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11206w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11211w11218w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11211w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11211w11214w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11211w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11076w11083w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11076w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11076w11079w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11076w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11216w11223w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11216w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11216w11219w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11216w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11221w11228w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11221w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11221w11224w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11221w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11226w11233w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11226w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11226w11229w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11226w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11231w11238w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11231w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11231w11234w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11231w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11236w11243w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11236w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11236w11239w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11236w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11241w11248w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11241w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11241w11244w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11241w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11246w11253w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11246w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11246w11249w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11246w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11251w11258w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11251w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11251w11254w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11251w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11256w11263w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11256w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11256w11259w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11256w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11261w11268w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11261w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11261w11264w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11261w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11081w11088w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11081w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11081w11084w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11081w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11266w11273w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11266w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11266w11269w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11266w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11271w11278w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11271w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11271w11274w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11271w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11276w11283w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11276w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11276w11279w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11276w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11281w11288w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11281w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11281w11284w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11281w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11286w11293w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11286w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11286w11289w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11286w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11291w11298w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11291w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11291w11294w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11291w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11296w11303w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11296w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11296w11299w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11296w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11301w11308w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11301w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11301w11304w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11301w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11306w11313w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11306w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11306w11309w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11306w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11311w11318w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11311w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11311w11314w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11311w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11086w11093w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11086w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11086w11089w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11086w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11316w11323w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11316w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11316w11319w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11316w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11321w11328w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11321w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11321w11324w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11321w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11326w11333w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11326w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11326w11329w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11326w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11331w11338w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11331w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11331w11334w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11331w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11336w11343w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11336w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11336w11339w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11336w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11341w11348w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11341w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11341w11344w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11341w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11346w11353w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11346w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11346w11349w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11346w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11351w11358w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11351w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11351w11354w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11351w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11356w11363w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11356w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11356w11359w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11356w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11361w11368w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11361w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11361w11364w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11361w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11091w11098w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11091w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11091w11094w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11091w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11366w11373w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11366w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11366w11369w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11366w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11371w11378w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11371w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11371w11374w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11371w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11376w11383w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11376w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11376w11379w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11376w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11381w11388w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11381w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11381w11384w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11381w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11386w11393w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11386w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11386w11389w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11386w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11391w11398w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11391w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11391w11394w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11391w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11396w11403w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11396w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11396w11399w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11396w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11401w11408w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11401w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11401w11404w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11401w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11406w11413w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11406w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11406w11409w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11406w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11411w11418w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11411w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11411w11414w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11411w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11096w11103w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11096w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11096w11099w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11096w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11416w11423w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11416w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11416w11419w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11416w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11421w11428w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11421w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11421w11424w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11421w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11426w11433w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11426w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11426w11429w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11426w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11431w11438w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11431w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11431w11434w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11431w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11436w11443w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11436w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11436w11439w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11436w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11441w11448w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11441w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11441w11444w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11441w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11446w11453w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11446w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11446w11449w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11446w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11451w11457w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11451w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11451w11454w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11451w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11458w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11048w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11101w11108w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11101w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11101w11104w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11101w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11106w11113w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11106w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11106w11109w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11106w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11111w11118w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11111w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11111w11114w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11111w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w(0) <= NOT wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w11120w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11116w11119w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11111w11118w(0);
	wire_crr_fp_range1_w11125w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11121w11124w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11116w11123w(0);
	wire_crr_fp_range1_w11130w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11126w11129w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11121w11128w(0);
	wire_crr_fp_range1_w11135w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11131w11134w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11126w11133w(0);
	wire_crr_fp_range1_w11140w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11136w11139w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11131w11138w(0);
	wire_crr_fp_range1_w11145w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11141w11144w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11136w11143w(0);
	wire_crr_fp_range1_w11150w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11146w11149w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11141w11148w(0);
	wire_crr_fp_range1_w11155w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11151w11154w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11146w11153w(0);
	wire_crr_fp_range1_w11160w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11156w11159w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11151w11158w(0);
	wire_crr_fp_range1_w11165w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11161w11164w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11156w11163w(0);
	wire_crr_fp_range1_w11074w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11070w11073w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11069w11072w(0);
	wire_crr_fp_range1_w11170w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11166w11169w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11161w11168w(0);
	wire_crr_fp_range1_w11175w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11171w11174w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11166w11173w(0);
	wire_crr_fp_range1_w11180w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11176w11179w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11171w11178w(0);
	wire_crr_fp_range1_w11185w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11181w11184w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11176w11183w(0);
	wire_crr_fp_range1_w11190w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11186w11189w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11181w11188w(0);
	wire_crr_fp_range1_w11195w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11191w11194w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11186w11193w(0);
	wire_crr_fp_range1_w11200w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11196w11199w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11191w11198w(0);
	wire_crr_fp_range1_w11205w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11201w11204w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11196w11203w(0);
	wire_crr_fp_range1_w11210w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11206w11209w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11201w11208w(0);
	wire_crr_fp_range1_w11215w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11211w11214w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11206w11213w(0);
	wire_crr_fp_range1_w11080w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11076w11079w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11070w11078w(0);
	wire_crr_fp_range1_w11220w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11216w11219w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11211w11218w(0);
	wire_crr_fp_range1_w11225w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11221w11224w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11216w11223w(0);
	wire_crr_fp_range1_w11230w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11226w11229w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11221w11228w(0);
	wire_crr_fp_range1_w11235w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11231w11234w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11226w11233w(0);
	wire_crr_fp_range1_w11240w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11236w11239w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11231w11238w(0);
	wire_crr_fp_range1_w11245w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11241w11244w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11236w11243w(0);
	wire_crr_fp_range1_w11250w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11246w11249w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11241w11248w(0);
	wire_crr_fp_range1_w11255w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11251w11254w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11246w11253w(0);
	wire_crr_fp_range1_w11260w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11256w11259w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11251w11258w(0);
	wire_crr_fp_range1_w11265w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11261w11264w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11256w11263w(0);
	wire_crr_fp_range1_w11085w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11081w11084w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11076w11083w(0);
	wire_crr_fp_range1_w11270w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11266w11269w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11261w11268w(0);
	wire_crr_fp_range1_w11275w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11271w11274w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11266w11273w(0);
	wire_crr_fp_range1_w11280w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11276w11279w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11271w11278w(0);
	wire_crr_fp_range1_w11285w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11281w11284w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11276w11283w(0);
	wire_crr_fp_range1_w11290w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11286w11289w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11281w11288w(0);
	wire_crr_fp_range1_w11295w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11291w11294w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11286w11293w(0);
	wire_crr_fp_range1_w11300w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11296w11299w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11291w11298w(0);
	wire_crr_fp_range1_w11305w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11301w11304w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11296w11303w(0);
	wire_crr_fp_range1_w11310w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11306w11309w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11301w11308w(0);
	wire_crr_fp_range1_w11315w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11311w11314w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11306w11313w(0);
	wire_crr_fp_range1_w11090w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11086w11089w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11081w11088w(0);
	wire_crr_fp_range1_w11320w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11316w11319w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11311w11318w(0);
	wire_crr_fp_range1_w11325w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11321w11324w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11316w11323w(0);
	wire_crr_fp_range1_w11330w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11326w11329w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11321w11328w(0);
	wire_crr_fp_range1_w11335w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11331w11334w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11326w11333w(0);
	wire_crr_fp_range1_w11340w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11336w11339w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11331w11338w(0);
	wire_crr_fp_range1_w11345w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11341w11344w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11336w11343w(0);
	wire_crr_fp_range1_w11350w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11346w11349w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11341w11348w(0);
	wire_crr_fp_range1_w11355w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11351w11354w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11346w11353w(0);
	wire_crr_fp_range1_w11360w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11356w11359w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11351w11358w(0);
	wire_crr_fp_range1_w11365w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11361w11364w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11356w11363w(0);
	wire_crr_fp_range1_w11095w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11091w11094w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11086w11093w(0);
	wire_crr_fp_range1_w11370w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11366w11369w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11361w11368w(0);
	wire_crr_fp_range1_w11375w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11371w11374w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11366w11373w(0);
	wire_crr_fp_range1_w11380w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11376w11379w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11371w11378w(0);
	wire_crr_fp_range1_w11385w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11381w11384w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11376w11383w(0);
	wire_crr_fp_range1_w11390w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11386w11389w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11381w11388w(0);
	wire_crr_fp_range1_w11395w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11391w11394w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11386w11393w(0);
	wire_crr_fp_range1_w11400w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11396w11399w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11391w11398w(0);
	wire_crr_fp_range1_w11405w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11401w11404w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11396w11403w(0);
	wire_crr_fp_range1_w11410w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11406w11409w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11401w11408w(0);
	wire_crr_fp_range1_w11415w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11411w11414w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11406w11413w(0);
	wire_crr_fp_range1_w11100w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11096w11099w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11091w11098w(0);
	wire_crr_fp_range1_w11420w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11416w11419w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11411w11418w(0);
	wire_crr_fp_range1_w11425w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11421w11424w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11416w11423w(0);
	wire_crr_fp_range1_w11430w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11426w11429w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11421w11428w(0);
	wire_crr_fp_range1_w11435w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11431w11434w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11426w11433w(0);
	wire_crr_fp_range1_w11440w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11436w11439w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11431w11438w(0);
	wire_crr_fp_range1_w11445w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11441w11444w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11436w11443w(0);
	wire_crr_fp_range1_w11450w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11446w11449w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11441w11448w(0);
	wire_crr_fp_range1_w11455w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11451w11454w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11446w11453w(0);
	wire_crr_fp_range1_w11459w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11458w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11451w11457w(0);
	wire_crr_fp_range1_w11105w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11101w11104w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11096w11103w(0);
	wire_crr_fp_range1_w11110w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11106w11109w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11101w11108w(0);
	wire_crr_fp_range1_w11115w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11111w11114w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11106w11113w(0);
	basefractiondelnode_w <= cbfd_5;
	basefractionnode_w <= wire_fp_range_table1_basefraction;
	circle <= circleff(35 DOWNTO 0);
	circlenode_w <= wire_circle_add_result;
	const_23_w <= "000010111";
	incexponentnode_w <= wire_fp_range_table1_incexponent;
	incmantissanode_w <= wire_fp_range_table1_incmantissa;
	leadnode_w <= (NOT wire_clz23_q);
	mantissaexponentnode_w <= wire_exponent_adjust_sub_result;
	mantissamultipliernode_w <= wire_csftin_result;
	multipliernode_w <= wire_mult23x56_result;
	multipliernormnode_w <= ( wire_crr_fp_range1_w11459w & wire_crr_fp_range1_w11455w & wire_crr_fp_range1_w11450w & wire_crr_fp_range1_w11445w & wire_crr_fp_range1_w11440w & wire_crr_fp_range1_w11435w & wire_crr_fp_range1_w11430w & wire_crr_fp_range1_w11425w & wire_crr_fp_range1_w11420w & wire_crr_fp_range1_w11415w & wire_crr_fp_range1_w11410w & wire_crr_fp_range1_w11405w & wire_crr_fp_range1_w11400w & wire_crr_fp_range1_w11395w & wire_crr_fp_range1_w11390w & wire_crr_fp_range1_w11385w & wire_crr_fp_range1_w11380w & wire_crr_fp_range1_w11375w & wire_crr_fp_range1_w11370w & wire_crr_fp_range1_w11365w & wire_crr_fp_range1_w11360w & wire_crr_fp_range1_w11355w & wire_crr_fp_range1_w11350w & wire_crr_fp_range1_w11345w & wire_crr_fp_range1_w11340w & wire_crr_fp_range1_w11335w & wire_crr_fp_range1_w11330w & wire_crr_fp_range1_w11325w & wire_crr_fp_range1_w11320w & wire_crr_fp_range1_w11315w & wire_crr_fp_range1_w11310w & wire_crr_fp_range1_w11305w & wire_crr_fp_range1_w11300w & wire_crr_fp_range1_w11295w & wire_crr_fp_range1_w11290w & wire_crr_fp_range1_w11285w & wire_crr_fp_range1_w11280w & wire_crr_fp_range1_w11275w & wire_crr_fp_range1_w11270w & wire_crr_fp_range1_w11265w & wire_crr_fp_range1_w11260w & wire_crr_fp_range1_w11255w & wire_crr_fp_range1_w11250w & wire_crr_fp_range1_w11245w & wire_crr_fp_range1_w11240w & wire_crr_fp_range1_w11235w & wire_crr_fp_range1_w11230w & wire_crr_fp_range1_w11225w & wire_crr_fp_range1_w11220w & wire_crr_fp_range1_w11215w & wire_crr_fp_range1_w11210w & wire_crr_fp_range1_w11205w & wire_crr_fp_range1_w11200w & wire_crr_fp_range1_w11195w & wire_crr_fp_range1_w11190w & wire_crr_fp_range1_w11185w & wire_crr_fp_range1_w11180w & wire_crr_fp_range1_w11175w & wire_crr_fp_range1_w11170w & wire_crr_fp_range1_w11165w & wire_crr_fp_range1_w11160w & wire_crr_fp_range1_w11155w & wire_crr_fp_range1_w11150w & wire_crr_fp_range1_w11145w & wire_crr_fp_range1_w11140w & wire_crr_fp_range1_w11135w & wire_crr_fp_range1_w11130w & wire_crr_fp_range1_w11125w & wire_crr_fp_range1_w11120w & wire_crr_fp_range1_w11115w
 & wire_crr_fp_range1_w11110w & wire_crr_fp_range1_w11105w & wire_crr_fp_range1_w11100w & wire_crr_fp_range1_w11095w & wire_crr_fp_range1_w11090w & wire_crr_fp_range1_w11085w & wire_crr_fp_range1_w11080w & wire_crr_fp_range1_w11074w);
	negbasefractiondelnode_w <= wire_negbasedractiondel_sub_result;
	negcircle <= negcircleff(35 DOWNTO 0);
	negcirclenode_w <= wire_negcircle_add_result;
	negrotatenode_w <= ( wire_rotateff_w_lg_w_q_range11583w11585w & wire_rotateff_w_lg_w_q_range11580w11582w & wire_rotateff_w_lg_w_q_range11577w11579w & wire_rotateff_w_lg_w_q_range11574w11576w & wire_rotateff_w_lg_w_q_range11571w11573w & wire_rotateff_w_lg_w_q_range11568w11570w & wire_rotateff_w_lg_w_q_range11565w11567w & wire_rotateff_w_lg_w_q_range11562w11564w & wire_rotateff_w_lg_w_q_range11559w11561w & wire_rotateff_w_lg_w_q_range11556w11558w & wire_rotateff_w_lg_w_q_range11553w11555w & wire_rotateff_w_lg_w_q_range11550w11552w & wire_rotateff_w_lg_w_q_range11547w11549w & wire_rotateff_w_lg_w_q_range11544w11546w & wire_rotateff_w_lg_w_q_range11541w11543w & wire_rotateff_w_lg_w_q_range11538w11540w & wire_rotateff_w_lg_w_q_range11535w11537w & wire_rotateff_w_lg_w_q_range11532w11534w & wire_rotateff_w_lg_w_q_range11529w11531w & wire_rotateff_w_lg_w_q_range11526w11528w & wire_rotateff_w_lg_w_q_range11523w11525w & wire_rotateff_w_lg_w_q_range11520w11522w & wire_rotateff_w_lg_w_q_range11517w11519w & wire_rotateff_w_lg_w_q_range11514w11516w & wire_rotateff_w_lg_w_q_range11511w11513w & wire_rotateff_w_lg_w_q_range11508w11510w & wire_rotateff_w_lg_w_q_range11505w11507w & wire_rotateff_w_lg_w_q_range11502w11504w & wire_rotateff_w_lg_w_q_range11499w11501w & wire_rotateff_w_lg_w_q_range11496w11498w & wire_rotateff_w_lg_w_q_range11493w11495w & wire_rotateff_w_lg_w_q_range11490w11492w & wire_rotateff_w_lg_w_q_range11487w11489w & wire_rotateff_w_lg_w_q_range11484w11486w & wire_rotateff_w_lg_w_q_range11481w11483w & wire_rotateff_w_lg_w_q_range11477w11479w);
	rotatenode_w <= wire_fp_lsft_rsft78_result;
	wire_crr_fp_range1_w_data_range11039w <= data(22 DOWNTO 0);
	wire_crr_fp_range1_w_data_range11040w <= data(30 DOWNTO 23);
	wire_crr_fp_range1_w_multipliernode_w_range11069w(0) <= multipliernode_w(0);
	wire_crr_fp_range1_w_multipliernode_w_range11116w(0) <= multipliernode_w(10);
	wire_crr_fp_range1_w_multipliernode_w_range11121w(0) <= multipliernode_w(11);
	wire_crr_fp_range1_w_multipliernode_w_range11126w(0) <= multipliernode_w(12);
	wire_crr_fp_range1_w_multipliernode_w_range11131w(0) <= multipliernode_w(13);
	wire_crr_fp_range1_w_multipliernode_w_range11136w(0) <= multipliernode_w(14);
	wire_crr_fp_range1_w_multipliernode_w_range11141w(0) <= multipliernode_w(15);
	wire_crr_fp_range1_w_multipliernode_w_range11146w(0) <= multipliernode_w(16);
	wire_crr_fp_range1_w_multipliernode_w_range11151w(0) <= multipliernode_w(17);
	wire_crr_fp_range1_w_multipliernode_w_range11156w(0) <= multipliernode_w(18);
	wire_crr_fp_range1_w_multipliernode_w_range11161w(0) <= multipliernode_w(19);
	wire_crr_fp_range1_w_multipliernode_w_range11070w(0) <= multipliernode_w(1);
	wire_crr_fp_range1_w_multipliernode_w_range11166w(0) <= multipliernode_w(20);
	wire_crr_fp_range1_w_multipliernode_w_range11171w(0) <= multipliernode_w(21);
	wire_crr_fp_range1_w_multipliernode_w_range11176w(0) <= multipliernode_w(22);
	wire_crr_fp_range1_w_multipliernode_w_range11181w(0) <= multipliernode_w(23);
	wire_crr_fp_range1_w_multipliernode_w_range11186w(0) <= multipliernode_w(24);
	wire_crr_fp_range1_w_multipliernode_w_range11191w(0) <= multipliernode_w(25);
	wire_crr_fp_range1_w_multipliernode_w_range11196w(0) <= multipliernode_w(26);
	wire_crr_fp_range1_w_multipliernode_w_range11201w(0) <= multipliernode_w(27);
	wire_crr_fp_range1_w_multipliernode_w_range11206w(0) <= multipliernode_w(28);
	wire_crr_fp_range1_w_multipliernode_w_range11211w(0) <= multipliernode_w(29);
	wire_crr_fp_range1_w_multipliernode_w_range11076w(0) <= multipliernode_w(2);
	wire_crr_fp_range1_w_multipliernode_w_range11216w(0) <= multipliernode_w(30);
	wire_crr_fp_range1_w_multipliernode_w_range11221w(0) <= multipliernode_w(31);
	wire_crr_fp_range1_w_multipliernode_w_range11226w(0) <= multipliernode_w(32);
	wire_crr_fp_range1_w_multipliernode_w_range11231w(0) <= multipliernode_w(33);
	wire_crr_fp_range1_w_multipliernode_w_range11236w(0) <= multipliernode_w(34);
	wire_crr_fp_range1_w_multipliernode_w_range11241w(0) <= multipliernode_w(35);
	wire_crr_fp_range1_w_multipliernode_w_range11246w(0) <= multipliernode_w(36);
	wire_crr_fp_range1_w_multipliernode_w_range11251w(0) <= multipliernode_w(37);
	wire_crr_fp_range1_w_multipliernode_w_range11256w(0) <= multipliernode_w(38);
	wire_crr_fp_range1_w_multipliernode_w_range11261w(0) <= multipliernode_w(39);
	wire_crr_fp_range1_w_multipliernode_w_range11081w(0) <= multipliernode_w(3);
	wire_crr_fp_range1_w_multipliernode_w_range11266w(0) <= multipliernode_w(40);
	wire_crr_fp_range1_w_multipliernode_w_range11271w(0) <= multipliernode_w(41);
	wire_crr_fp_range1_w_multipliernode_w_range11276w(0) <= multipliernode_w(42);
	wire_crr_fp_range1_w_multipliernode_w_range11281w(0) <= multipliernode_w(43);
	wire_crr_fp_range1_w_multipliernode_w_range11286w(0) <= multipliernode_w(44);
	wire_crr_fp_range1_w_multipliernode_w_range11291w(0) <= multipliernode_w(45);
	wire_crr_fp_range1_w_multipliernode_w_range11296w(0) <= multipliernode_w(46);
	wire_crr_fp_range1_w_multipliernode_w_range11301w(0) <= multipliernode_w(47);
	wire_crr_fp_range1_w_multipliernode_w_range11306w(0) <= multipliernode_w(48);
	wire_crr_fp_range1_w_multipliernode_w_range11311w(0) <= multipliernode_w(49);
	wire_crr_fp_range1_w_multipliernode_w_range11086w(0) <= multipliernode_w(4);
	wire_crr_fp_range1_w_multipliernode_w_range11316w(0) <= multipliernode_w(50);
	wire_crr_fp_range1_w_multipliernode_w_range11321w(0) <= multipliernode_w(51);
	wire_crr_fp_range1_w_multipliernode_w_range11326w(0) <= multipliernode_w(52);
	wire_crr_fp_range1_w_multipliernode_w_range11331w(0) <= multipliernode_w(53);
	wire_crr_fp_range1_w_multipliernode_w_range11336w(0) <= multipliernode_w(54);
	wire_crr_fp_range1_w_multipliernode_w_range11341w(0) <= multipliernode_w(55);
	wire_crr_fp_range1_w_multipliernode_w_range11346w(0) <= multipliernode_w(56);
	wire_crr_fp_range1_w_multipliernode_w_range11351w(0) <= multipliernode_w(57);
	wire_crr_fp_range1_w_multipliernode_w_range11356w(0) <= multipliernode_w(58);
	wire_crr_fp_range1_w_multipliernode_w_range11361w(0) <= multipliernode_w(59);
	wire_crr_fp_range1_w_multipliernode_w_range11091w(0) <= multipliernode_w(5);
	wire_crr_fp_range1_w_multipliernode_w_range11366w(0) <= multipliernode_w(60);
	wire_crr_fp_range1_w_multipliernode_w_range11371w(0) <= multipliernode_w(61);
	wire_crr_fp_range1_w_multipliernode_w_range11376w(0) <= multipliernode_w(62);
	wire_crr_fp_range1_w_multipliernode_w_range11381w(0) <= multipliernode_w(63);
	wire_crr_fp_range1_w_multipliernode_w_range11386w(0) <= multipliernode_w(64);
	wire_crr_fp_range1_w_multipliernode_w_range11391w(0) <= multipliernode_w(65);
	wire_crr_fp_range1_w_multipliernode_w_range11396w(0) <= multipliernode_w(66);
	wire_crr_fp_range1_w_multipliernode_w_range11401w(0) <= multipliernode_w(67);
	wire_crr_fp_range1_w_multipliernode_w_range11406w(0) <= multipliernode_w(68);
	wire_crr_fp_range1_w_multipliernode_w_range11411w(0) <= multipliernode_w(69);
	wire_crr_fp_range1_w_multipliernode_w_range11096w(0) <= multipliernode_w(6);
	wire_crr_fp_range1_w_multipliernode_w_range11416w(0) <= multipliernode_w(70);
	wire_crr_fp_range1_w_multipliernode_w_range11421w(0) <= multipliernode_w(71);
	wire_crr_fp_range1_w_multipliernode_w_range11426w(0) <= multipliernode_w(72);
	wire_crr_fp_range1_w_multipliernode_w_range11431w(0) <= multipliernode_w(73);
	wire_crr_fp_range1_w_multipliernode_w_range11436w(0) <= multipliernode_w(74);
	wire_crr_fp_range1_w_multipliernode_w_range11441w(0) <= multipliernode_w(75);
	wire_crr_fp_range1_w_multipliernode_w_range11446w(0) <= multipliernode_w(76);
	wire_crr_fp_range1_w_multipliernode_w_range11451w(0) <= multipliernode_w(77);
	wire_crr_fp_range1_w_multipliernode_w_range11048w(0) <= multipliernode_w(78);
	wire_crr_fp_range1_w_multipliernode_w_range11101w(0) <= multipliernode_w(7);
	wire_crr_fp_range1_w_multipliernode_w_range11106w(0) <= multipliernode_w(8);
	wire_crr_fp_range1_w_multipliernode_w_range11111w(0) <= multipliernode_w(9);
	fp_range_table1 :  mysincos_altfp_sincos_srrt_gra
	  PORT MAP ( 
		address => tableaddressff,
		basefraction => wire_fp_range_table1_basefraction,
		incexponent => wire_fp_range_table1_incexponent,
		incmantissa => wire_fp_range_table1_incmantissa
	  );
	wire_clz23_data <= ( mantissaff & "111111111");
	clz23 :  mysincos_altpriority_encoder_qb6
	  PORT MAP ( 
		data => wire_clz23_data,
		q => wire_clz23_q
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN basefractiondelff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN basefractiondelff <= basefractiondelnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN basefractionff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN basefractionff <= basefractionnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cbfd_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cbfd_0 <= basefractionff;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cbfd_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cbfd_1 <= cbfd_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cbfd_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cbfd_2 <= cbfd_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cbfd_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cbfd_3 <= cbfd_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cbfd_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cbfd_4 <= cbfd_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cbfd_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cbfd_5 <= cbfd_4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN circleff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN circleff <= circlenode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponentff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN exponentff <= wire_crr_fp_range1_w_data_range11040w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN incexponentff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN incexponentff <= incexponentnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN incmantissaff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN incmantissaff <= incmantissanode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN leadff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN leadff <= leadnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissadelff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN mantissadelff <= mantissaff;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissaff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN mantissaff <= wire_crr_fp_range1_w_data_range11039w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissamultiplierff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN mantissamultiplierff <= mantissamultipliernode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN multipliernormff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN multipliernormff <= multipliernormnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN negbasefractiondelff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN negbasefractiondelff <= negbasefractiondelnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN negcircleff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN negcircleff <= negcirclenode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN negrangeexponentff4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN negrangeexponentff4 <= wire_negrangeexponent_sub4_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN negrangeexponentff5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN negrangeexponentff5 <= wire_negrangeexponent_sub5_result;
			END IF;
		END IF;
	END PROCESS;
	loop53 : FOR i IN 0 TO 6 GENERATE 
		wire_negrangeexponentff5_w_lg_w_lg_w_q_range11460w11464w11465w(i) <= wire_negrangeexponentff5_w_lg_w_q_range11460w11464w(0) AND wire_rangeexponentff_5_w_q_range11463w(i);
	END GENERATE loop53;
	loop54 : FOR i IN 0 TO 6 GENERATE 
		wire_negrangeexponentff5_w_lg_w_q_range11460w11462w(i) <= wire_negrangeexponentff5_w_q_range11460w(0) AND wire_negrangeexponentff5_w_q_range11461w(i);
	END GENERATE loop54;
	wire_negrangeexponentff5_w_lg_w_q_range11460w11464w(0) <= NOT wire_negrangeexponentff5_w_q_range11460w(0);
	wire_negrangeexponentff5_w_q_range11461w <= negrangeexponentff5(6 DOWNTO 0);
	wire_negrangeexponentff5_w_q_range11460w(0) <= negrangeexponentff5(8);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rangeexponentff_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rangeexponentff_0 <= mantissaexponentnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rangeexponentff_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rangeexponentff_1 <= wire_rangeexponent_sub1_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rangeexponentff_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rangeexponentff_2 <= rangeexponentff_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rangeexponentff_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rangeexponentff_3 <= rangeexponentff_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rangeexponentff_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rangeexponentff_4 <= rangeexponentff_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rangeexponentff_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rangeexponentff_5 <= wire_rangeexponent_sub5_result;
			END IF;
		END IF;
	END PROCESS;
	wire_rangeexponentff_5_w_q_range11463w <= rangeexponentff_5(6 DOWNTO 0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rotateff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rotateff <= rotatenode_w;
			END IF;
		END IF;
	END PROCESS;
	wire_rotateff_w_lg_w_q_range11477w11479w(0) <= NOT wire_rotateff_w_q_range11477w(0);
	wire_rotateff_w_lg_w_q_range11481w11483w(0) <= NOT wire_rotateff_w_q_range11481w(0);
	wire_rotateff_w_lg_w_q_range11484w11486w(0) <= NOT wire_rotateff_w_q_range11484w(0);
	wire_rotateff_w_lg_w_q_range11487w11489w(0) <= NOT wire_rotateff_w_q_range11487w(0);
	wire_rotateff_w_lg_w_q_range11490w11492w(0) <= NOT wire_rotateff_w_q_range11490w(0);
	wire_rotateff_w_lg_w_q_range11493w11495w(0) <= NOT wire_rotateff_w_q_range11493w(0);
	wire_rotateff_w_lg_w_q_range11496w11498w(0) <= NOT wire_rotateff_w_q_range11496w(0);
	wire_rotateff_w_lg_w_q_range11499w11501w(0) <= NOT wire_rotateff_w_q_range11499w(0);
	wire_rotateff_w_lg_w_q_range11502w11504w(0) <= NOT wire_rotateff_w_q_range11502w(0);
	wire_rotateff_w_lg_w_q_range11505w11507w(0) <= NOT wire_rotateff_w_q_range11505w(0);
	wire_rotateff_w_lg_w_q_range11508w11510w(0) <= NOT wire_rotateff_w_q_range11508w(0);
	wire_rotateff_w_lg_w_q_range11511w11513w(0) <= NOT wire_rotateff_w_q_range11511w(0);
	wire_rotateff_w_lg_w_q_range11514w11516w(0) <= NOT wire_rotateff_w_q_range11514w(0);
	wire_rotateff_w_lg_w_q_range11517w11519w(0) <= NOT wire_rotateff_w_q_range11517w(0);
	wire_rotateff_w_lg_w_q_range11520w11522w(0) <= NOT wire_rotateff_w_q_range11520w(0);
	wire_rotateff_w_lg_w_q_range11523w11525w(0) <= NOT wire_rotateff_w_q_range11523w(0);
	wire_rotateff_w_lg_w_q_range11526w11528w(0) <= NOT wire_rotateff_w_q_range11526w(0);
	wire_rotateff_w_lg_w_q_range11529w11531w(0) <= NOT wire_rotateff_w_q_range11529w(0);
	wire_rotateff_w_lg_w_q_range11532w11534w(0) <= NOT wire_rotateff_w_q_range11532w(0);
	wire_rotateff_w_lg_w_q_range11535w11537w(0) <= NOT wire_rotateff_w_q_range11535w(0);
	wire_rotateff_w_lg_w_q_range11538w11540w(0) <= NOT wire_rotateff_w_q_range11538w(0);
	wire_rotateff_w_lg_w_q_range11541w11543w(0) <= NOT wire_rotateff_w_q_range11541w(0);
	wire_rotateff_w_lg_w_q_range11544w11546w(0) <= NOT wire_rotateff_w_q_range11544w(0);
	wire_rotateff_w_lg_w_q_range11547w11549w(0) <= NOT wire_rotateff_w_q_range11547w(0);
	wire_rotateff_w_lg_w_q_range11550w11552w(0) <= NOT wire_rotateff_w_q_range11550w(0);
	wire_rotateff_w_lg_w_q_range11553w11555w(0) <= NOT wire_rotateff_w_q_range11553w(0);
	wire_rotateff_w_lg_w_q_range11556w11558w(0) <= NOT wire_rotateff_w_q_range11556w(0);
	wire_rotateff_w_lg_w_q_range11559w11561w(0) <= NOT wire_rotateff_w_q_range11559w(0);
	wire_rotateff_w_lg_w_q_range11562w11564w(0) <= NOT wire_rotateff_w_q_range11562w(0);
	wire_rotateff_w_lg_w_q_range11565w11567w(0) <= NOT wire_rotateff_w_q_range11565w(0);
	wire_rotateff_w_lg_w_q_range11568w11570w(0) <= NOT wire_rotateff_w_q_range11568w(0);
	wire_rotateff_w_lg_w_q_range11571w11573w(0) <= NOT wire_rotateff_w_q_range11571w(0);
	wire_rotateff_w_lg_w_q_range11574w11576w(0) <= NOT wire_rotateff_w_q_range11574w(0);
	wire_rotateff_w_lg_w_q_range11577w11579w(0) <= NOT wire_rotateff_w_q_range11577w(0);
	wire_rotateff_w_lg_w_q_range11580w11582w(0) <= NOT wire_rotateff_w_q_range11580w(0);
	wire_rotateff_w_lg_w_q_range11583w11585w(0) <= NOT wire_rotateff_w_q_range11583w(0);
	wire_rotateff_w_q_range11477w(0) <= rotateff(42);
	wire_rotateff_w_q_range11481w(0) <= rotateff(43);
	wire_rotateff_w_q_range11484w(0) <= rotateff(44);
	wire_rotateff_w_q_range11487w(0) <= rotateff(45);
	wire_rotateff_w_q_range11490w(0) <= rotateff(46);
	wire_rotateff_w_q_range11493w(0) <= rotateff(47);
	wire_rotateff_w_q_range11496w(0) <= rotateff(48);
	wire_rotateff_w_q_range11499w(0) <= rotateff(49);
	wire_rotateff_w_q_range11502w(0) <= rotateff(50);
	wire_rotateff_w_q_range11505w(0) <= rotateff(51);
	wire_rotateff_w_q_range11508w(0) <= rotateff(52);
	wire_rotateff_w_q_range11511w(0) <= rotateff(53);
	wire_rotateff_w_q_range11514w(0) <= rotateff(54);
	wire_rotateff_w_q_range11517w(0) <= rotateff(55);
	wire_rotateff_w_q_range11520w(0) <= rotateff(56);
	wire_rotateff_w_q_range11523w(0) <= rotateff(57);
	wire_rotateff_w_q_range11526w(0) <= rotateff(58);
	wire_rotateff_w_q_range11529w(0) <= rotateff(59);
	wire_rotateff_w_q_range11532w(0) <= rotateff(60);
	wire_rotateff_w_q_range11535w(0) <= rotateff(61);
	wire_rotateff_w_q_range11538w(0) <= rotateff(62);
	wire_rotateff_w_q_range11541w(0) <= rotateff(63);
	wire_rotateff_w_q_range11544w(0) <= rotateff(64);
	wire_rotateff_w_q_range11547w(0) <= rotateff(65);
	wire_rotateff_w_q_range11550w(0) <= rotateff(66);
	wire_rotateff_w_q_range11553w(0) <= rotateff(67);
	wire_rotateff_w_q_range11556w(0) <= rotateff(68);
	wire_rotateff_w_q_range11559w(0) <= rotateff(69);
	wire_rotateff_w_q_range11562w(0) <= rotateff(70);
	wire_rotateff_w_q_range11565w(0) <= rotateff(71);
	wire_rotateff_w_q_range11568w(0) <= rotateff(72);
	wire_rotateff_w_q_range11571w(0) <= rotateff(73);
	wire_rotateff_w_q_range11574w(0) <= rotateff(74);
	wire_rotateff_w_q_range11577w(0) <= rotateff(75);
	wire_rotateff_w_q_range11580w(0) <= rotateff(76);
	wire_rotateff_w_q_range11583w(0) <= rotateff(77);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN tableaddressff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN tableaddressff <= exponentff;
			END IF;
		END IF;
	END PROCESS;
	wire_circle_add_dataa <= ( "0" & basefractiondelff);
	wire_circle_add_datab <= ( "0" & rotateff(77 DOWNTO 42));
	circle_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 37
	  )
	  PORT MAP ( 
		dataa => wire_circle_add_dataa,
		datab => wire_circle_add_datab,
		result => wire_circle_add_result
	  );
	wire_exponent_adjust_sub_datab <= ( "0000" & leadff);
	exponent_adjust_sub :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => const_23_w,
		datab => wire_exponent_adjust_sub_datab,
		result => wire_exponent_adjust_sub_result
	  );
	wire_negbasedractiondel_sub_dataa <= (OTHERS => '0');
	negbasedractiondel_sub :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 36
	  )
	  PORT MAP ( 
		dataa => wire_negbasedractiondel_sub_dataa,
		datab => basefractiondelnode_w(35 DOWNTO 0),
		result => wire_negbasedractiondel_sub_result
	  );
	wire_negcircle_add_dataa <= ( "1" & negbasefractiondelff);
	wire_negcircle_add_datab <= ( "1" & negrotatenode_w);
	negcircle_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 37
	  )
	  PORT MAP ( 
		cin => wire_vcc,
		dataa => wire_negcircle_add_dataa,
		datab => wire_negcircle_add_datab,
		result => wire_negcircle_add_result
	  );
	wire_negrangeexponent_sub4_dataa <= ( "1" & "00000000");
	negrangeexponent_sub4 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => wire_negrangeexponent_sub4_dataa,
		datab => rangeexponentff_3,
		result => wire_negrangeexponent_sub4_result
	  );
	wire_negrangeexponent_sub5_datab <= ( "00000000" & wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w);
	negrangeexponent_sub5 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => negrangeexponentff4,
		datab => wire_negrangeexponent_sub5_datab,
		result => wire_negrangeexponent_sub5_result
	  );
	wire_rangeexponent_sub1_datab <= ( "0" & incexponentff);
	rangeexponent_sub1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => rangeexponentff_0,
		datab => wire_rangeexponent_sub1_datab,
		result => wire_rangeexponent_sub1_result
	  );
	wire_rangeexponent_sub5_datab <= ( "00000000" & wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11050w);
	rangeexponent_sub5 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => rangeexponentff_4,
		datab => wire_rangeexponent_sub5_datab,
		result => wire_rangeexponent_sub5_result
	  );
	csftin :  lpm_clshift
	  GENERIC MAP (
		LPM_WIDTH => 23,
		LPM_WIDTHDIST => 5
	  )
	  PORT MAP ( 
		data => mantissadelff,
		direction => wire_gnd,
		distance => leadff,
		result => wire_csftin_result
	  );
	wire_fp_lsft_rsft78_distance <= wire_negrangeexponentff5_w_lg_w_lg_w_lg_w_q_range11460w11464w11465w11466w;
	loop55 : FOR i IN 0 TO 6 GENERATE 
		wire_negrangeexponentff5_w_lg_w_lg_w_lg_w_q_range11460w11464w11465w11466w(i) <= wire_negrangeexponentff5_w_lg_w_lg_w_q_range11460w11464w11465w(i) OR wire_negrangeexponentff5_w_lg_w_q_range11460w11462w(i);
	END GENERATE loop55;
	fp_lsft_rsft78 :  lpm_clshift
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_WIDTH => 78,
		LPM_WIDTHDIST => 7
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		data => multipliernormff,
		direction => negrangeexponentff5(8),
		distance => wire_fp_lsft_rsft78_distance,
		result => wire_fp_lsft_rsft78_result
	  );
	mult23x56 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 4,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 23,
		LPM_WIDTHB => 56,
		LPM_WIDTHP => 79
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => mantissamultiplierff,
		datab => incmantissaff,
		result => wire_mult23x56_result
	  );

 END RTL; --mysincos_altfp_sincos_range_79c


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" WIDTH=64 WIDTHAD=6 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=32 WIDTHAD=5 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altpriority_encoder_q08 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0)
	 ); 
 END mysincos_altpriority_encoder_q08;

 ARCHITECTURE RTL OF mysincos_altpriority_encoder_q08 IS

	 SIGNAL  wire_altpriority_encoder19_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_w_lg_zero13074w13075w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_zero13076w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_zero13074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_w_lg_zero13076w13077w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_zero	:	STD_LOGIC;
	 COMPONENT  mysincos_altpriority_encoder_r08
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  mysincos_altpriority_encoder_rf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder20_w_lg_zero13074w & wire_altpriority_encoder20_w_lg_w_lg_zero13076w13077w);
	altpriority_encoder19 :  mysincos_altpriority_encoder_r08
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder19_q
	  );
	loop56 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder20_w_lg_w_lg_zero13074w13075w(i) <= wire_altpriority_encoder20_w_lg_zero13074w(0) AND wire_altpriority_encoder20_q(i);
	END GENERATE loop56;
	loop57 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder20_w_lg_zero13076w(i) <= wire_altpriority_encoder20_zero AND wire_altpriority_encoder19_q(i);
	END GENERATE loop57;
	wire_altpriority_encoder20_w_lg_zero13074w(0) <= NOT wire_altpriority_encoder20_zero;
	loop58 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder20_w_lg_w_lg_zero13076w13077w(i) <= wire_altpriority_encoder20_w_lg_zero13076w(i) OR wire_altpriority_encoder20_w_lg_w_lg_zero13074w13075w(i);
	END GENERATE loop58;
	altpriority_encoder20 :  mysincos_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder20_q,
		zero => wire_altpriority_encoder20_zero
	  );

 END RTL; --mysincos_altpriority_encoder_q08


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=32 WIDTHAD=5 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altpriority_encoder_qf8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END mysincos_altpriority_encoder_qf8;

 ARCHITECTURE RTL OF mysincos_altpriority_encoder_qf8 IS

	 SIGNAL  wire_altpriority_encoder21_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder21_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder22_w_lg_w_lg_zero13083w13084w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_zero13085w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_zero13083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_w_lg_zero13085w13086w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_zero	:	STD_LOGIC;
	 COMPONENT  mysincos_altpriority_encoder_rf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder22_w_lg_zero13083w & wire_altpriority_encoder22_w_lg_w_lg_zero13085w13086w);
	zero <= (wire_altpriority_encoder21_zero AND wire_altpriority_encoder22_zero);
	altpriority_encoder21 :  mysincos_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder21_q,
		zero => wire_altpriority_encoder21_zero
	  );
	loop59 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder22_w_lg_w_lg_zero13083w13084w(i) <= wire_altpriority_encoder22_w_lg_zero13083w(0) AND wire_altpriority_encoder22_q(i);
	END GENERATE loop59;
	loop60 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder22_w_lg_zero13085w(i) <= wire_altpriority_encoder22_zero AND wire_altpriority_encoder21_q(i);
	END GENERATE loop60;
	wire_altpriority_encoder22_w_lg_zero13083w(0) <= NOT wire_altpriority_encoder22_zero;
	loop61 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder22_w_lg_w_lg_zero13085w13086w(i) <= wire_altpriority_encoder22_w_lg_zero13085w(i) OR wire_altpriority_encoder22_w_lg_w_lg_zero13083w13084w(i);
	END GENERATE loop61;
	altpriority_encoder22 :  mysincos_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder22_q,
		zero => wire_altpriority_encoder22_zero
	  );

 END RTL; --mysincos_altpriority_encoder_qf8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altpriority_encoder_0c6 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (63 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (5 DOWNTO 0)
	 ); 
 END mysincos_altpriority_encoder_0c6;

 ARCHITECTURE RTL OF mysincos_altpriority_encoder_0c6 IS

	 SIGNAL  wire_altpriority_encoder17_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_w_lg_zero13065w13066w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_zero13067w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_zero13065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_w_lg_zero13067w13068w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_zero	:	STD_LOGIC;
	 COMPONENT  mysincos_altpriority_encoder_q08
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  mysincos_altpriority_encoder_qf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder18_w_lg_zero13065w & wire_altpriority_encoder18_w_lg_w_lg_zero13067w13068w);
	altpriority_encoder17 :  mysincos_altpriority_encoder_q08
	  PORT MAP ( 
		data => data(31 DOWNTO 0),
		q => wire_altpriority_encoder17_q
	  );
	loop62 : FOR i IN 0 TO 4 GENERATE 
		wire_altpriority_encoder18_w_lg_w_lg_zero13065w13066w(i) <= wire_altpriority_encoder18_w_lg_zero13065w(0) AND wire_altpriority_encoder18_q(i);
	END GENERATE loop62;
	loop63 : FOR i IN 0 TO 4 GENERATE 
		wire_altpriority_encoder18_w_lg_zero13067w(i) <= wire_altpriority_encoder18_zero AND wire_altpriority_encoder17_q(i);
	END GENERATE loop63;
	wire_altpriority_encoder18_w_lg_zero13065w(0) <= NOT wire_altpriority_encoder18_zero;
	loop64 : FOR i IN 0 TO 4 GENERATE 
		wire_altpriority_encoder18_w_lg_w_lg_zero13067w13068w(i) <= wire_altpriority_encoder18_w_lg_zero13067w(i) OR wire_altpriority_encoder18_w_lg_w_lg_zero13065w13066w(i);
	END GENERATE loop64;
	altpriority_encoder18 :  mysincos_altpriority_encoder_qf8
	  PORT MAP ( 
		data => data(63 DOWNTO 32),
		q => wire_altpriority_encoder18_q,
		zero => wire_altpriority_encoder18_zero
	  );

 END RTL; --mysincos_altpriority_encoder_0c6

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 52 lpm_clshift 3 lpm_mult 3 lpm_mux 2 reg 3720 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  mysincos_altfp_sincos_0ae IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END mysincos_altfp_sincos_0ae;

 ARCHITECTURE RTL OF mysincos_altfp_sincos_0ae IS

	 SIGNAL  wire_ccc_cordic_m_sincos	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_circle	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_negcircle	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_clz_data	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_clz_q	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL	 countff	:	STD_LOGIC_VECTOR(5 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exponentinff	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exponentnormff	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exponentnormff_w_lg_q398w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_exponentnormff_w_lg_w_lg_q398w399w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 exponentoutff	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 fixed_sincosff	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_0	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_1	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_10	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_11	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_12	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_13	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_14	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_15	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_16	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_17	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_18	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_19	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_2	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_20	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_21	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_22	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_23	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_24	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_25	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_26	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_27	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_28	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_29	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_3	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_30	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_31	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_32	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_33	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_34	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_4	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_5	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_6	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_7	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_8	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_9	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mantissanormff	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_mantissanormff_w_lg_q394w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_mantissanormff_w_lg_w_lg_q394w395w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL	 mantissaoutff	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 quadrant_sumff	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 select_sincosff	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 selectoutputff	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_selectoutputff_w_lg_w_q_range390w393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_selectoutputff_w_q_range390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 signcalcff	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_signcalcff_w_lg_w_q_range401w403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_signcalcff_w_q_range401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 signinff	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_signinff_w_q_range56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 signoutff	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exponentcheck_sub_dataa	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_exponentcheck_sub_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_exponentcheck_sub_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_exponentnorm_add_datab	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_exponentnorm_add_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_exponentnormmode_sub_datab	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_exponentnormmode_sub_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_mantissanorm_add_datab	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_mantissanorm_add_result	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_quadrantsum_add_cin	:	STD_LOGIC;
	 SIGNAL  wire_quadrantsum_add_result	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_sft_result	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_cmul_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_w_lg_negative_quadrant_w19w	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_w_lg_positive_quadrant_w20w	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_circle_w_range7w8w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_input_number_delay_w_range391w392w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_input_number_delay_w_range396w397w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range311w313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range314w316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range317w319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range320w322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range323w325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range326w328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range329w331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range332w334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range335w337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range338w340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range341w343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range344w346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range347w349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range350w352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range353w355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range356w358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range359w361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range362w364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range365w367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range368w370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range371w373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range374w376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range377w379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_negcircle_w_range4w5w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_w_lg_quadrantselect_w6w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_quadrant_w_range17w18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range249w252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range278w282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range281w285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range284w288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range287w291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range290w294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range251w255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range254w258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range257w261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range260w264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range263w267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range266w270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range269w273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range272w276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range275w279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_quadrantsign_w58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  aclr	:	STD_LOGIC;
	 SIGNAL  circle_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  countnode_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  exponentcheck_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exponentnormmode_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  fixed_sincos_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  fixed_sincosnode_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  fraction_quadrant_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  indexbit_w :	STD_LOGIC;
	 SIGNAL  indexcheck_w :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  input_number_delay_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  input_number_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  mantissanormnode_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  negative_quadrant_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  negcircle_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  one_term_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  overflownode_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  piovertwo_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  positive_quadrant_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  quadrant_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  quadrantselect_w :	STD_LOGIC;
	 SIGNAL  quadrantsign_w :	STD_LOGIC;
	 SIGNAL  radiansnode_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  value_128_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  value_x73_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  zerovec_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_w_circle_w_range7w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_w_data_range128w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_input_number_delay_w_range391w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_input_number_delay_w_range396w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_negcircle_w_range4w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_quadrant_w_range17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  mysincos_altfp_sincos_cordic_m_a8e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		indexbit	:	IN  STD_LOGIC := '0';
		radians	:	IN  STD_LOGIC_VECTOR(33 DOWNTO 0) := (OTHERS => '0');
		sincos	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		sincosbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  mysincos_altfp_sincos_range_79c
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		circle	:	OUT  STD_LOGIC_VECTOR(35 DOWNTO 0);
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
		negcircle	:	OUT  STD_LOGIC_VECTOR(35 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  mysincos_altpriority_encoder_0c6
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(63 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(5 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_clshift
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_SHIFTTYPE	:	STRING := "LOGICAL";
		LPM_WIDTH	:	NATURAL;
		LPM_WIDTHDIST	:	NATURAL;
		lpm_type	:	STRING := "lpm_clshift"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		direction	:	IN STD_LOGIC := '0';
		distance	:	IN STD_LOGIC_VECTOR(LPM_WIDTHDIST-1 DOWNTO 0);
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		underflow	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_mult
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTHA	:	NATURAL;
		LPM_WIDTHB	:	NATURAL;
		LPM_WIDTHP	:	NATURAL;
		LPM_WIDTHS	:	NATURAL := 1;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_mult"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTHA-1 DOWNTO 0);
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTHB-1 DOWNTO 0);
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHP-1 DOWNTO 0);
		sum	:	IN STD_LOGIC_VECTOR(LPM_WIDTHS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	loop65 : FOR i IN 0 TO 35 GENERATE 
		wire_w_lg_negative_quadrant_w19w(i) <= negative_quadrant_w(i) AND wire_w_lg_w_quadrant_w_range17w18w(0);
	END GENERATE loop65;
	loop66 : FOR i IN 0 TO 35 GENERATE 
		wire_w_lg_positive_quadrant_w20w(i) <= positive_quadrant_w(i) AND wire_w_quadrant_w_range17w(0);
	END GENERATE loop66;
	loop67 : FOR i IN 0 TO 33 GENERATE 
		wire_w_lg_w_circle_w_range7w8w(i) <= wire_w_circle_w_range7w(i) AND wire_w_lg_quadrantselect_w6w(0);
	END GENERATE loop67;
	loop68 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_w_input_number_delay_w_range391w392w(i) <= wire_w_input_number_delay_w_range391w(i) AND wire_selectoutputff_w_q_range390w(0);
	END GENERATE loop68;
	loop69 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_input_number_delay_w_range396w397w(i) <= wire_w_input_number_delay_w_range396w(i) AND wire_selectoutputff_w_q_range390w(0);
	END GENERATE loop69;
	wire_w_lg_w_mantissanormnode_w_range311w313w(0) <= wire_w_mantissanormnode_w_range311w(0) AND wire_w_overflownode_w_range309w(0);
	wire_w_lg_w_mantissanormnode_w_range314w316w(0) <= wire_w_mantissanormnode_w_range314w(0) AND wire_w_overflownode_w_range312w(0);
	wire_w_lg_w_mantissanormnode_w_range317w319w(0) <= wire_w_mantissanormnode_w_range317w(0) AND wire_w_overflownode_w_range315w(0);
	wire_w_lg_w_mantissanormnode_w_range320w322w(0) <= wire_w_mantissanormnode_w_range320w(0) AND wire_w_overflownode_w_range318w(0);
	wire_w_lg_w_mantissanormnode_w_range323w325w(0) <= wire_w_mantissanormnode_w_range323w(0) AND wire_w_overflownode_w_range321w(0);
	wire_w_lg_w_mantissanormnode_w_range326w328w(0) <= wire_w_mantissanormnode_w_range326w(0) AND wire_w_overflownode_w_range324w(0);
	wire_w_lg_w_mantissanormnode_w_range329w331w(0) <= wire_w_mantissanormnode_w_range329w(0) AND wire_w_overflownode_w_range327w(0);
	wire_w_lg_w_mantissanormnode_w_range332w334w(0) <= wire_w_mantissanormnode_w_range332w(0) AND wire_w_overflownode_w_range330w(0);
	wire_w_lg_w_mantissanormnode_w_range335w337w(0) <= wire_w_mantissanormnode_w_range335w(0) AND wire_w_overflownode_w_range333w(0);
	wire_w_lg_w_mantissanormnode_w_range338w340w(0) <= wire_w_mantissanormnode_w_range338w(0) AND wire_w_overflownode_w_range336w(0);
	wire_w_lg_w_mantissanormnode_w_range341w343w(0) <= wire_w_mantissanormnode_w_range341w(0) AND wire_w_overflownode_w_range339w(0);
	wire_w_lg_w_mantissanormnode_w_range344w346w(0) <= wire_w_mantissanormnode_w_range344w(0) AND wire_w_overflownode_w_range342w(0);
	wire_w_lg_w_mantissanormnode_w_range347w349w(0) <= wire_w_mantissanormnode_w_range347w(0) AND wire_w_overflownode_w_range345w(0);
	wire_w_lg_w_mantissanormnode_w_range350w352w(0) <= wire_w_mantissanormnode_w_range350w(0) AND wire_w_overflownode_w_range348w(0);
	wire_w_lg_w_mantissanormnode_w_range353w355w(0) <= wire_w_mantissanormnode_w_range353w(0) AND wire_w_overflownode_w_range351w(0);
	wire_w_lg_w_mantissanormnode_w_range356w358w(0) <= wire_w_mantissanormnode_w_range356w(0) AND wire_w_overflownode_w_range354w(0);
	wire_w_lg_w_mantissanormnode_w_range359w361w(0) <= wire_w_mantissanormnode_w_range359w(0) AND wire_w_overflownode_w_range357w(0);
	wire_w_lg_w_mantissanormnode_w_range362w364w(0) <= wire_w_mantissanormnode_w_range362w(0) AND wire_w_overflownode_w_range360w(0);
	wire_w_lg_w_mantissanormnode_w_range365w367w(0) <= wire_w_mantissanormnode_w_range365w(0) AND wire_w_overflownode_w_range363w(0);
	wire_w_lg_w_mantissanormnode_w_range368w370w(0) <= wire_w_mantissanormnode_w_range368w(0) AND wire_w_overflownode_w_range366w(0);
	wire_w_lg_w_mantissanormnode_w_range371w373w(0) <= wire_w_mantissanormnode_w_range371w(0) AND wire_w_overflownode_w_range369w(0);
	wire_w_lg_w_mantissanormnode_w_range374w376w(0) <= wire_w_mantissanormnode_w_range374w(0) AND wire_w_overflownode_w_range372w(0);
	wire_w_lg_w_mantissanormnode_w_range377w379w(0) <= wire_w_mantissanormnode_w_range377w(0) AND wire_w_overflownode_w_range375w(0);
	loop70 : FOR i IN 0 TO 33 GENERATE 
		wire_w_lg_w_negcircle_w_range4w5w(i) <= wire_w_negcircle_w_range4w(i) AND quadrantselect_w;
	END GENERATE loop70;
	wire_w_lg_quadrantselect_w6w(0) <= NOT quadrantselect_w;
	wire_w_lg_w_quadrant_w_range17w18w(0) <= NOT wire_w_quadrant_w_range17w(0);
	wire_w_lg_w_indexcheck_w_range249w252w(0) <= wire_w_indexcheck_w_range249w(0) OR wire_w_radiansnode_w_range248w(0);
	wire_w_lg_w_indexcheck_w_range278w282w(0) <= wire_w_indexcheck_w_range278w(0) OR wire_w_radiansnode_w_range280w(0);
	wire_w_lg_w_indexcheck_w_range281w285w(0) <= wire_w_indexcheck_w_range281w(0) OR wire_w_radiansnode_w_range283w(0);
	wire_w_lg_w_indexcheck_w_range284w288w(0) <= wire_w_indexcheck_w_range284w(0) OR wire_w_radiansnode_w_range286w(0);
	wire_w_lg_w_indexcheck_w_range287w291w(0) <= wire_w_indexcheck_w_range287w(0) OR wire_w_radiansnode_w_range289w(0);
	wire_w_lg_w_indexcheck_w_range290w294w(0) <= wire_w_indexcheck_w_range290w(0) OR wire_w_radiansnode_w_range292w(0);
	wire_w_lg_w_indexcheck_w_range251w255w(0) <= wire_w_indexcheck_w_range251w(0) OR wire_w_radiansnode_w_range253w(0);
	wire_w_lg_w_indexcheck_w_range254w258w(0) <= wire_w_indexcheck_w_range254w(0) OR wire_w_radiansnode_w_range256w(0);
	wire_w_lg_w_indexcheck_w_range257w261w(0) <= wire_w_indexcheck_w_range257w(0) OR wire_w_radiansnode_w_range259w(0);
	wire_w_lg_w_indexcheck_w_range260w264w(0) <= wire_w_indexcheck_w_range260w(0) OR wire_w_radiansnode_w_range262w(0);
	wire_w_lg_w_indexcheck_w_range263w267w(0) <= wire_w_indexcheck_w_range263w(0) OR wire_w_radiansnode_w_range265w(0);
	wire_w_lg_w_indexcheck_w_range266w270w(0) <= wire_w_indexcheck_w_range266w(0) OR wire_w_radiansnode_w_range268w(0);
	wire_w_lg_w_indexcheck_w_range269w273w(0) <= wire_w_indexcheck_w_range269w(0) OR wire_w_radiansnode_w_range271w(0);
	wire_w_lg_w_indexcheck_w_range272w276w(0) <= wire_w_indexcheck_w_range272w(0) OR wire_w_radiansnode_w_range274w(0);
	wire_w_lg_w_indexcheck_w_range275w279w(0) <= wire_w_indexcheck_w_range275w(0) OR wire_w_radiansnode_w_range277w(0);
	wire_w_lg_quadrantsign_w58w(0) <= quadrantsign_w XOR wire_signinff_w_q_range56w(0);
	aclr <= '0';
	circle_w <= wire_crr_fp_range1_circle;
	clk_en <= '1';
	countnode_w <= (NOT wire_clz_q);
	exponentcheck_w <= wire_exponentcheck_sub_result;
	exponentnormmode_w <= wire_exponentnormmode_sub_result;
	fixed_sincos_w <= wire_ccc_cordic_m_sincos;
	fixed_sincosnode_w <= ( fixed_sincos_w & zerovec_w(1 DOWNTO 0));
	fraction_quadrant_w <= (wire_w_lg_positive_quadrant_w20w OR wire_w_lg_negative_quadrant_w19w);
	indexbit_w <= (NOT indexcheck_w(3));
	indexcheck_w <= ( wire_w_lg_w_indexcheck_w_range290w294w & wire_w_lg_w_indexcheck_w_range287w291w & wire_w_lg_w_indexcheck_w_range284w288w & wire_w_lg_w_indexcheck_w_range281w285w & wire_w_lg_w_indexcheck_w_range278w282w & wire_w_lg_w_indexcheck_w_range275w279w & wire_w_lg_w_indexcheck_w_range272w276w & wire_w_lg_w_indexcheck_w_range269w273w & wire_w_lg_w_indexcheck_w_range266w270w & wire_w_lg_w_indexcheck_w_range263w267w & wire_w_lg_w_indexcheck_w_range260w264w & wire_w_lg_w_indexcheck_w_range257w261w & wire_w_lg_w_indexcheck_w_range254w258w & wire_w_lg_w_indexcheck_w_range251w255w & wire_w_lg_w_indexcheck_w_range249w252w & radiansnode_w(32));
	input_number_delay_w <= input_delay_ff_34;
	input_number_w <= data;
	mantissanormnode_w <= wire_sft_result;
	negative_quadrant_w <= (NOT positive_quadrant_w);
	negcircle_w <= wire_crr_fp_range1_negcircle;
	one_term_w <= ( wire_w_lg_w_quadrant_w_range17w18w & zerovec_w(34 DOWNTO 0));
	overflownode_w <= ( wire_w_lg_w_mantissanormnode_w_range377w379w & wire_w_lg_w_mantissanormnode_w_range374w376w & wire_w_lg_w_mantissanormnode_w_range371w373w & wire_w_lg_w_mantissanormnode_w_range368w370w & wire_w_lg_w_mantissanormnode_w_range365w367w & wire_w_lg_w_mantissanormnode_w_range362w364w & wire_w_lg_w_mantissanormnode_w_range359w361w & wire_w_lg_w_mantissanormnode_w_range356w358w & wire_w_lg_w_mantissanormnode_w_range353w355w & wire_w_lg_w_mantissanormnode_w_range350w352w & wire_w_lg_w_mantissanormnode_w_range347w349w & wire_w_lg_w_mantissanormnode_w_range344w346w & wire_w_lg_w_mantissanormnode_w_range341w343w & wire_w_lg_w_mantissanormnode_w_range338w340w & wire_w_lg_w_mantissanormnode_w_range335w337w & wire_w_lg_w_mantissanormnode_w_range332w334w & wire_w_lg_w_mantissanormnode_w_range329w331w & wire_w_lg_w_mantissanormnode_w_range326w328w & wire_w_lg_w_mantissanormnode_w_range323w325w & wire_w_lg_w_mantissanormnode_w_range320w322w & wire_w_lg_w_mantissanormnode_w_range317w319w & wire_w_lg_w_mantissanormnode_w_range314w316w & wire_w_lg_w_mantissanormnode_w_range311w313w & mantissanormnode_w(11));
	piovertwo_w <= "110010010000111111011010101000100010";
	positive_quadrant_w <= ( "0" & quadrant_w & "0");
	quadrant_w <= (wire_w_lg_w_circle_w_range7w8w OR wire_w_lg_w_negcircle_w_range4w5w);
	quadrantselect_w <= circle_w(34);
	quadrantsign_w <= circle_w(35);
	radiansnode_w <= wire_cmul_result;
	result <= ( signoutff & exponentoutff & mantissaoutff);
	value_128_w <= "10000000";
	value_x73_w <= "01110011";
	zerovec_w <= (OTHERS => '0');
	wire_w_circle_w_range7w <= circle_w(33 DOWNTO 0);
	wire_w_data_range128w <= data(30 DOWNTO 23);
	wire_w_indexcheck_w_range249w(0) <= indexcheck_w(0);
	wire_w_indexcheck_w_range278w(0) <= indexcheck_w(10);
	wire_w_indexcheck_w_range281w(0) <= indexcheck_w(11);
	wire_w_indexcheck_w_range284w(0) <= indexcheck_w(12);
	wire_w_indexcheck_w_range287w(0) <= indexcheck_w(13);
	wire_w_indexcheck_w_range290w(0) <= indexcheck_w(14);
	wire_w_indexcheck_w_range251w(0) <= indexcheck_w(1);
	wire_w_indexcheck_w_range254w(0) <= indexcheck_w(2);
	wire_w_indexcheck_w_range257w(0) <= indexcheck_w(3);
	wire_w_indexcheck_w_range260w(0) <= indexcheck_w(4);
	wire_w_indexcheck_w_range263w(0) <= indexcheck_w(5);
	wire_w_indexcheck_w_range266w(0) <= indexcheck_w(6);
	wire_w_indexcheck_w_range269w(0) <= indexcheck_w(7);
	wire_w_indexcheck_w_range272w(0) <= indexcheck_w(8);
	wire_w_indexcheck_w_range275w(0) <= indexcheck_w(9);
	wire_w_input_number_delay_w_range391w <= input_number_delay_w(22 DOWNTO 0);
	wire_w_input_number_delay_w_range396w <= input_number_delay_w(30 DOWNTO 23);
	wire_w_mantissanormnode_w_range311w(0) <= mantissanormnode_w(12);
	wire_w_mantissanormnode_w_range314w(0) <= mantissanormnode_w(13);
	wire_w_mantissanormnode_w_range317w(0) <= mantissanormnode_w(14);
	wire_w_mantissanormnode_w_range320w(0) <= mantissanormnode_w(15);
	wire_w_mantissanormnode_w_range323w(0) <= mantissanormnode_w(16);
	wire_w_mantissanormnode_w_range326w(0) <= mantissanormnode_w(17);
	wire_w_mantissanormnode_w_range329w(0) <= mantissanormnode_w(18);
	wire_w_mantissanormnode_w_range332w(0) <= mantissanormnode_w(19);
	wire_w_mantissanormnode_w_range335w(0) <= mantissanormnode_w(20);
	wire_w_mantissanormnode_w_range338w(0) <= mantissanormnode_w(21);
	wire_w_mantissanormnode_w_range341w(0) <= mantissanormnode_w(22);
	wire_w_mantissanormnode_w_range344w(0) <= mantissanormnode_w(23);
	wire_w_mantissanormnode_w_range347w(0) <= mantissanormnode_w(24);
	wire_w_mantissanormnode_w_range350w(0) <= mantissanormnode_w(25);
	wire_w_mantissanormnode_w_range353w(0) <= mantissanormnode_w(26);
	wire_w_mantissanormnode_w_range356w(0) <= mantissanormnode_w(27);
	wire_w_mantissanormnode_w_range359w(0) <= mantissanormnode_w(28);
	wire_w_mantissanormnode_w_range362w(0) <= mantissanormnode_w(29);
	wire_w_mantissanormnode_w_range365w(0) <= mantissanormnode_w(30);
	wire_w_mantissanormnode_w_range368w(0) <= mantissanormnode_w(31);
	wire_w_mantissanormnode_w_range371w(0) <= mantissanormnode_w(32);
	wire_w_mantissanormnode_w_range374w(0) <= mantissanormnode_w(33);
	wire_w_mantissanormnode_w_range377w(0) <= mantissanormnode_w(34);
	wire_w_negcircle_w_range4w <= negcircle_w(33 DOWNTO 0);
	wire_w_overflownode_w_range309w(0) <= overflownode_w(0);
	wire_w_overflownode_w_range339w(0) <= overflownode_w(10);
	wire_w_overflownode_w_range342w(0) <= overflownode_w(11);
	wire_w_overflownode_w_range345w(0) <= overflownode_w(12);
	wire_w_overflownode_w_range348w(0) <= overflownode_w(13);
	wire_w_overflownode_w_range351w(0) <= overflownode_w(14);
	wire_w_overflownode_w_range354w(0) <= overflownode_w(15);
	wire_w_overflownode_w_range357w(0) <= overflownode_w(16);
	wire_w_overflownode_w_range360w(0) <= overflownode_w(17);
	wire_w_overflownode_w_range363w(0) <= overflownode_w(18);
	wire_w_overflownode_w_range366w(0) <= overflownode_w(19);
	wire_w_overflownode_w_range312w(0) <= overflownode_w(1);
	wire_w_overflownode_w_range369w(0) <= overflownode_w(20);
	wire_w_overflownode_w_range372w(0) <= overflownode_w(21);
	wire_w_overflownode_w_range375w(0) <= overflownode_w(22);
	wire_w_overflownode_w_range315w(0) <= overflownode_w(2);
	wire_w_overflownode_w_range318w(0) <= overflownode_w(3);
	wire_w_overflownode_w_range321w(0) <= overflownode_w(4);
	wire_w_overflownode_w_range324w(0) <= overflownode_w(5);
	wire_w_overflownode_w_range327w(0) <= overflownode_w(6);
	wire_w_overflownode_w_range330w(0) <= overflownode_w(7);
	wire_w_overflownode_w_range333w(0) <= overflownode_w(8);
	wire_w_overflownode_w_range336w(0) <= overflownode_w(9);
	wire_w_quadrant_w_range17w(0) <= quadrant_w(33);
	wire_w_radiansnode_w_range292w(0) <= radiansnode_w(18);
	wire_w_radiansnode_w_range289w(0) <= radiansnode_w(19);
	wire_w_radiansnode_w_range286w(0) <= radiansnode_w(20);
	wire_w_radiansnode_w_range283w(0) <= radiansnode_w(21);
	wire_w_radiansnode_w_range280w(0) <= radiansnode_w(22);
	wire_w_radiansnode_w_range277w(0) <= radiansnode_w(23);
	wire_w_radiansnode_w_range274w(0) <= radiansnode_w(24);
	wire_w_radiansnode_w_range271w(0) <= radiansnode_w(25);
	wire_w_radiansnode_w_range268w(0) <= radiansnode_w(26);
	wire_w_radiansnode_w_range265w(0) <= radiansnode_w(27);
	wire_w_radiansnode_w_range262w(0) <= radiansnode_w(28);
	wire_w_radiansnode_w_range259w(0) <= radiansnode_w(29);
	wire_w_radiansnode_w_range256w(0) <= radiansnode_w(30);
	wire_w_radiansnode_w_range253w(0) <= radiansnode_w(31);
	wire_w_radiansnode_w_range248w(0) <= radiansnode_w(32);
	ccc_cordic_m :  mysincos_altfp_sincos_cordic_m_a8e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		indexbit => indexbit_w,
		radians => radiansnode_w,
		sincos => wire_ccc_cordic_m_sincos,
		sincosbit => select_sincosff(3)
	  );
	crr_fp_range1 :  mysincos_altfp_sincos_range_79c
	  PORT MAP ( 
		aclr => aclr,
		circle => wire_crr_fp_range1_circle,
		clken => clk_en,
		clock => clock,
		data => data,
		negcircle => wire_crr_fp_range1_negcircle
	  );
	wire_clz_data <= ( fixed_sincosnode_w & "1111111111111111111111111111");
	clz :  mysincos_altpriority_encoder_0c6
	  PORT MAP ( 
		data => wire_clz_data,
		q => wire_clz_q
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN countff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN countff <= countnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponentinff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponentinff <= wire_w_data_range128w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponentnormff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponentnormff <= wire_exponentnorm_add_result;
			END IF;
		END IF;
	END PROCESS;
	loop71 : FOR i IN 0 TO 7 GENERATE 
		wire_exponentnormff_w_lg_q398w(i) <= exponentnormff(i) AND wire_selectoutputff_w_lg_w_q_range390w393w(0);
	END GENERATE loop71;
	loop72 : FOR i IN 0 TO 7 GENERATE 
		wire_exponentnormff_w_lg_w_lg_q398w399w(i) <= wire_exponentnormff_w_lg_q398w(i) OR wire_w_lg_w_input_number_delay_w_range396w397w(i);
	END GENERATE loop72;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponentoutff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponentoutff <= wire_exponentnormff_w_lg_w_lg_q398w399w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN fixed_sincosff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN fixed_sincosff <= fixed_sincosnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_0 <= input_number_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_1 <= input_delay_ff_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_10 <= input_delay_ff_9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_11 <= input_delay_ff_10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_12 <= input_delay_ff_11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_13 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_13 <= input_delay_ff_12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_14 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_14 <= input_delay_ff_13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_15 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_15 <= input_delay_ff_14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_16 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_16 <= input_delay_ff_15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_17 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_17 <= input_delay_ff_16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_18 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_18 <= input_delay_ff_17;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_19 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_19 <= input_delay_ff_18;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_2 <= input_delay_ff_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_20 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_20 <= input_delay_ff_19;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_21 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_21 <= input_delay_ff_20;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_22 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_22 <= input_delay_ff_21;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_23 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_23 <= input_delay_ff_22;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_24 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_24 <= input_delay_ff_23;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_25 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_25 <= input_delay_ff_24;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_26 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_26 <= input_delay_ff_25;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_27 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_27 <= input_delay_ff_26;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_28 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_28 <= input_delay_ff_27;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_29 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_29 <= input_delay_ff_28;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_3 <= input_delay_ff_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_30 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_30 <= input_delay_ff_29;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_31 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_31 <= input_delay_ff_30;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_32 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_32 <= input_delay_ff_31;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_33 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_33 <= input_delay_ff_32;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_34 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_34 <= input_delay_ff_33;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_4 <= input_delay_ff_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_5 <= input_delay_ff_4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_6 <= input_delay_ff_5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_7 <= input_delay_ff_6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_8 <= input_delay_ff_7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_9 <= input_delay_ff_8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissanormff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mantissanormff <= wire_mantissanorm_add_result;
			END IF;
		END IF;
	END PROCESS;
	loop73 : FOR i IN 0 TO 22 GENERATE 
		wire_mantissanormff_w_lg_q394w(i) <= mantissanormff(i) AND wire_selectoutputff_w_lg_w_q_range390w393w(0);
	END GENERATE loop73;
	loop74 : FOR i IN 0 TO 22 GENERATE 
		wire_mantissanormff_w_lg_w_lg_q394w395w(i) <= wire_mantissanormff_w_lg_q394w(i) OR wire_w_lg_w_input_number_delay_w_range391w392w(i);
	END GENERATE loop74;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissaoutff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mantissaoutff <= wire_mantissanormff_w_lg_w_lg_q394w395w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN quadrant_sumff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN quadrant_sumff <= wire_quadrantsum_add_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN select_sincosff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN select_sincosff <= ( select_sincosff(2 DOWNTO 0) & quadrant_w(33));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN selectoutputff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN selectoutputff <= ( selectoutputff(32 DOWNTO 0) & exponentcheck_w(8));
			END IF;
		END IF;
	END PROCESS;
	wire_selectoutputff_w_lg_w_q_range390w393w(0) <= NOT wire_selectoutputff_w_q_range390w(0);
	wire_selectoutputff_w_q_range390w(0) <= selectoutputff(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN signcalcff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN signcalcff <= ( signcalcff(22 DOWNTO 0) & wire_w_lg_quadrantsign_w58w);
			END IF;
		END IF;
	END PROCESS;
	wire_signcalcff_w_lg_w_q_range401w403w(0) <= wire_signcalcff_w_q_range401w(0) AND wire_selectoutputff_w_lg_w_q_range390w393w(0);
	wire_signcalcff_w_q_range401w(0) <= signcalcff(23);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN signinff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN signinff <= ( signinff(9 DOWNTO 0) & data(31));
			END IF;
		END IF;
	END PROCESS;
	wire_signinff_w_q_range56w(0) <= signinff(10);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN signoutff <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN signoutff <= (wire_signcalcff_w_lg_w_q_range401w403w(0) OR (input_number_delay_w(31) AND selectoutputff(33)));
			END IF;
		END IF;
	END PROCESS;
	wire_exponentcheck_sub_dataa <= ( "0" & exponentinff);
	wire_exponentcheck_sub_datab <= ( "0" & value_x73_w);
	exponentcheck_sub :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => wire_exponentcheck_sub_dataa,
		datab => wire_exponentcheck_sub_datab,
		result => wire_exponentcheck_sub_result
	  );
	wire_exponentnorm_add_datab <= ( "0000000" & overflownode_w(23));
	exponentnorm_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		dataa => exponentnormmode_w(7 DOWNTO 0),
		datab => wire_exponentnorm_add_datab,
		result => wire_exponentnorm_add_result
	  );
	wire_exponentnormmode_sub_datab <= ( "00" & countff);
	exponentnormmode_sub :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		dataa => value_128_w,
		datab => wire_exponentnormmode_sub_datab,
		result => wire_exponentnormmode_sub_result
	  );
	wire_mantissanorm_add_datab <= ( "0000000000000000000000" & mantissanormnode_w(11));
	mantissanorm_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 23
	  )
	  PORT MAP ( 
		dataa => mantissanormnode_w(34 DOWNTO 12),
		datab => wire_mantissanorm_add_datab,
		result => wire_mantissanorm_add_result
	  );
	wire_quadrantsum_add_cin <= wire_w_lg_w_quadrant_w_range17w18w(0);
	quadrantsum_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 36
	  )
	  PORT MAP ( 
		cin => wire_quadrantsum_add_cin,
		dataa => one_term_w,
		datab => fraction_quadrant_w,
		result => wire_quadrantsum_add_result
	  );
	sft :  lpm_clshift
	  GENERIC MAP (
		LPM_WIDTH => 36,
		LPM_WIDTHDIST => 6
	  )
	  PORT MAP ( 
		data => fixed_sincosff,
		direction => wire_gnd,
		distance => countff,
		result => wire_sft_result
	  );
	cmul :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 3,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 36,
		LPM_WIDTHB => 36,
		LPM_WIDTHP => 34
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => quadrant_sumff,
		datab => piovertwo_w,
		result => wire_cmul_result
	  );

 END RTL; --mysincos_altfp_sincos_0ae
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY mysincos IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		data		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END mysincos;


ARCHITECTURE RTL OF mysincos IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);



	COMPONENT mysincos_altfp_sincos_0ae
	PORT (
			clock	: IN STD_LOGIC ;
			data	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(31 DOWNTO 0);

	mysincos_altfp_sincos_0ae_component : mysincos_altfp_sincos_0ae
	PORT MAP (
		clock => clock,
		data => data,
		result => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: FPM_FORMAT NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: CONSTANT: OPERATION STRING "SIN"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "36"
-- Retrieval info: CONSTANT: ROUNDING STRING "TO_NEAREST"
-- Retrieval info: CONSTANT: WIDTH_EXP NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_MAN NUMERIC "23"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: data 0 0 32 0 INPUT NODEFVAL "data[31..0]"
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @data 0 0 32 0 data 0 0 32 0
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL mysincos.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mysincos.inc TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mysincos.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mysincos.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mysincos_inst.vhd TRUE
-- Retrieval info: LIB_FILE: lpm
