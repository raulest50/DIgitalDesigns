myclk_inst : myclk PORT MAP (
		ena	 => ena_sig,
		inclk	 => inclk_sig,
		outclk	 => outclk_sig
	);
